LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY SHIFT_LEFT1 IS 
    PORT (
        IN_SIGNAL : IN STD_LOGIC_VECTOR(12 DOWNTO 0);
        OUT_SIGNAL : OUT STD_LOGIC_VECTOR(14 DOWNTO 0)
    );
END SHIFT_LEFT2;

ARCHITECTURE Behavior OF SHIFT_LEFT2 IS

SIGNAL AUX1 : STD_LOGIC; 

BEGIN
    
    OUT_SIGNAL <= IN_SIGNAL(12 downto 0) & "0";

END Behavior;
