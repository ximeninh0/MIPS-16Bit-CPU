LIBRARY ieee;
use ieee.std_logic_1164.all;

PACKAGE CONSTANTS_PACKAGE IS

constant WORD_SIZE     : integer := 16;
constant ADDR_SIZE     : integer := 4;
constant BYTE_SIZE     : integer := 8;
CONSTANT INSTRUCT_QTD  : integer := 14;
END CONSTANTS_PACKAGE;
