LIBRARY ieee;
USE ieee.std_logic_1164.all;
use work.CPU_PACKAGE.all;

ENTITY REG_BANK IS 
	port(
			REG_READ1,REG_READ2 :IN STD_LOGIC_VECTOR(1 DOWNTO 0);
			WRITE_REG :IN STD_LOGIC_VECTOR(1 DOWNTO 0);
			WRITE_DATA :IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			REG_WRITE,REG_READ: IN STD_LOGIC;
			DATA_READ1 :OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
			DATA_READ2 :OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END REG_BANK;

ARCHITECTURE Behavior OF REG_BANK IS
SIGNAL R_IN,WRITE_AUX: STD_LOGIC_VECTOR(1 TO 3);
SIGNAL R1,R2,R3 : STD_LOGIC_VECTOR(3 DOWNTO 0);
BEGIN

	WITH WRITE_REG SELECT
		WRITE_AUX <= 	"001" WHEN "01",
							"010" WHEN "10",
							"100" WHEN "11",
							"000" WHEN OTHERS;

	
	R_IN(1) <= WRITE_AUX(1) AND REG_WRITE;
	R_IN(2) <= WRITE_AUX(2) AND REG_WRITE;
	R_IN(3) <= WRITE_AUX(3) AND REG_WRITE;

	REG1_INSTANCE: REG PORT MAP(WRITE_DATA,R_in(1),RESET,CLOCK,R1);
	REG2_INSTANCE: REG PORT MAP(WRITE_DATA,R_in(2),RESET,CLOCK,R2);
	REG3_INSTANCE: REG PORT MAP(WRITE_DATA,R_in(3),RESET,CLOCK,R3);

	WITH REG_READ1 SELECT
	 MUX1 <= R1 when "01",
				R2 when "10",
				R3 when "11",
				"000" when others;

	WITH REG_READ2 SELECT
	 MUX2 <= R1 when "01",
				R2 when "10",
				R3 when "11",
				"000" when others;
							
	BUFFER1_INSTANCE: BUFFER_TRI PORT MAP(MUX1,REG_READ,DATA_READ1);
	BUFFER2_INSTANCE: BUFFER_TRI PORT MAP(MUX2,REG_READ,DATA_READ2);

END Behavior;
