LIBRARY ieee;
USE ieee.std_logic_1164.all;
use work.CPU_PACKAGE.all;

ENTITY HAZARD_DETECTION_UNIT IS 
    port(
--			INSTRUCTION : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
			ID_EX_MEM_READ : IN STD_LOGIC;
			ID_EX_RT 	: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
			IF_ID_RS 	: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
			IF_ID_RT 	: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
			
			BUBBLE 		: OUT STD_LOGIC;
			PC_WRITE 	: OUT STD_LOGIC;
			IF_ID_WRITE : OUT STD_LOGIC
    );
END HAZARD_DETECTION_UNIT;


ARCHITECTURE Behavior OF HAZARD_DETECTION_UNIT IS
BEGIN
--    PC_WRITE <= '1';    
--    IF_ID_WRITE <= '1';
--	 BUBBLE <='0';
	 
	PROCESS(ALL)
	BEGIN
	IF (ID_EX_MEM_READ = '1' AND ((ID_EX_RT = IF_ID_RS) OR (ID_EX_RT = IF_ID_RT))) THEN
		PC_WRITE <= '0';
		IF_ID_WRITE <= '0';
		BUBBLE <= '1';
	ELSE
	    PC_WRITE <= '1';    
		 IF_ID_WRITE <= '1';
		 BUBBLE <='0';
	END IF;
	END PROCESS;

END Behavior;
