LIBRARY ieee;
USE ieee.std_logic_1164.all;
use work.CPU_PACKAGE.all;

ENTITY HAZARD_DETECTION_UNIT IS 
    port(
			OPCODE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
			ID_EX_MEM_READ : IN STD_LOGIC;
			ID_EX_RT 	: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
			IF_ID_RS 	: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
			IF_ID_RT 	: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
			
		  REG_DST_EX_MEM : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		  REG_DST_MEM_WB : IN STD_LOGIC_VECTOR(3 DOWNTO 0);

		  WRITE_REG_EX_MEM : IN STD_LOGIC;
		  WRITE_REG_MEM_WB : IN STD_LOGIC;
			
			BUBBLE 		: OUT STD_LOGIC;
			PC_WRITE 	: OUT STD_LOGIC;
			IF_ID_WRITE : OUT STD_LOGIC
    );
END HAZARD_DETECTION_UNIT;


ARCHITECTURE Behavior OF HAZARD_DETECTION_UNIT IS
BEGIN
--    PC_WRITE <= '1';    
--    IF_ID_WRITE <= '1';
--	 BUBBLE <='0';
	 
	PROCESS(ALL)
	BEGIN
	IF (ID_EX_MEM_READ = '1' AND ((ID_EX_RT = IF_ID_RS) OR (ID_EX_RT = IF_ID_RT))) THEN
		PC_WRITE <= '0';
		IF_ID_WRITE <= '0';
		BUBBLE <= '1';
	ELSIF (WRITE_REG_EX_MEM = '1') AND (REG_DST_EX_MEM /= "0000") AND (REG_DST_EX_MEM = IF_ID_RS) AND OPCODE="100" THEN
			PC_WRITE <= '0';
		IF_ID_WRITE <= '0';
		BUBBLE <= '1';
	
	ELSIF (WRITE_REG_EX_MEM = '1') AND (REG_DST_EX_MEM /= "0000") AND (REG_DST_EX_MEM = IF_ID_RT) AND OPCODE="100" THEN
			PC_WRITE <= '0';
		IF_ID_WRITE <= '0';
		BUBBLE <= '1';
	ELSIF (WRITE_REG_MEM_WB = '1') AND (REG_DST_MEM_WB /= "0000") AND (REG_DST_MEM_WB = IF_ID_RS) AND OPCODE="100" THEN
			PC_WRITE <= '0';
		IF_ID_WRITE <= '0';
		BUBBLE <= '1';
	
	ELSIF (WRITE_REG_MEM_WB = '1') AND (REG_DST_MEM_WB /= "0000") AND (REG_DST_MEM_WB = IF_ID_RT) AND OPCODE="100" THEN
		PC_WRITE <= '0';
		IF_ID_WRITE <= '0';
		BUBBLE <= '1';
	ELSE
	    PC_WRITE <= '1';    
		 IF_ID_WRITE <= '1';
		 BUBBLE <='0';
	END IF;
	END PROCESS;

END Behavior;
