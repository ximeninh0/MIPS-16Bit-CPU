LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY CONTRACT_SIGNAL IS 
    PORT (
        IN_SIGNAL : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
        OUT_SIGNAL : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
    );
END CONTRACT_SIGNAL;

ARCHITECTURE Behavior OF CONTRACT_SIGNAL IS
BEGIN

    OUT_SIGNAL<= IN_SIGNAL(7 downto 0);

END Behavior;
