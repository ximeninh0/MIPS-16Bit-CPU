LIBRARY ieee;
use ieee.std_logic_1164.all;
use work.CONSTANTS_PACKAGE.all;
--PACKAGE COM TODOS OS COMPONENTES UTILIZADOS NA CPU E NA ULA

PACKAGE CPU_PACKAGE IS
	COMPONENT ULA IS 
		port(
				A,B : IN STD_LOGIC_VECTOR(15 DOWNTO 0);		-- Entradas A e B de 8 bits
				RESULT: out STD_LOGIC_VECTOR(15 DOWNTO 0);	-- Resultado de 4 bits
				OPERATION: IN STD_LOGIC;					-- Entrada que indica a operação que será realizada pela ULA
				ZERO, OVERFLOW,Cout : OUT STD_LOGIC		-- ZERO: 1 em caso do resultado ser 0, OV: 1 no caso da operação resultar em Overflow, Cout: 1 em caso de carry-out
			);
	END COMPONENT;
	
	COMPONENT UC_CPU IS 
		port(
			OPCODE : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			Clock : in std_logic;
			RESET : IN STD_LOGIC;
			En : IN STD_LOGIC;
			R_in : OUT STD_LOGIC_VECTOR(1 TO 3);
			R_out : OUT STD_LOGIC_VECTOR(1 TO 3);
			G_in : OUT STD_LOGIC;
			G_out : OUT STD_LOGIC;
			A_in : OUT STD_LOGIC;
			B_in : OUT STD_LOGIC;
			DONE : OUT STD_LOGIC;
			EXTERN : OUT STD_LOGIC;
			OP_ULA: OUT STD_LOGIC_VECTOR (3 DOWNTO 0)
		);
	END COMPONENT;
	
	COMPONENT UC_LCD IS 
		  port(
			OPCODE : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			 CLOCK : IN STD_LOGIC;
			 EQU,GRT,LST,ENABLE : IN STD_LOGIC;
			 LCD_DATA : out STD_LOGIC_VECTOR(7 DOWNTO 0);
			 LCD_RW : OUT STD_LOGIC;
			 LCD_EN : OUT STD_LOGIC;
			 LCD_RS: OUT STD_LOGIC
		  );
	END COMPONENT;
	
	COMPONENT AND_COMPONENT IS 
		port(
			X,Y :IN STD_LOGIC_VECTOR(15 DOWNTO 0);
			Z : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
		);
	END COMPONENT;
	
	COMPONENT OR_COMPONENT IS
		port(
			X,Y :IN STD_LOGIC_VECTOR(15 DOWNTO 0);
			Z : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
		);
	END COMPONENT;
	
	COMPONENT NOT_COMPONENT IS
		port(
			X,Y :IN STD_LOGIC_VECTOR(15 DOWNTO 0);
			Z : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
		);
	END COMPONENT;
	
	COMPONENT MULTI_COMPONENT IS
		port(
			X,Y :IN STD_LOGIC_VECTOR(1 DOWNTO 0);
			Z : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
		);
	END COMPONENT;
	
	
	COMPONENT RIPPLE_CARRY IS 
		port(
			A,B : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
			Cin : IN STD_LOGIC;
			Add_sub: IN STD_LOGIC;
			Overflow: OUT STD_LOGIC;
			Cout : OUT STD_LOGIC;
			Z : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
		);
	END COMPONENT;
	
	COMPONENT FULLADDER IS 
		port(
			A,B,Cin : IN STD_LOGIC;
			S,Cout : OUT STD_LOGIC
		);
	END COMPONENT;
	
	COMPONENT COMPARATOR16 IS 
		 port(
			  A,B : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
			  EQU : OUT STD_LOGIC
		 );
	END COMPONENT;
	
	COMPONENT SEGS_3_TRANSLATOR IS
		port(
			NUMBER : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
			TRANSLATED : OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
		);
	END COMPONENT;
	
	COMPONENT SEGS_4_TRANSLATOR IS 
		port(
			NUMBER : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
			TRANSLATED : OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
		);
	END COMPONENT;
	
	COMPONENT MUX_2_TO_1 IS 
		port(
			KEY : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
			X1,X2 : IN STD_LOGIC;
			F : OUT STD_LOGIC
		);
	END COMPONENT;
	
	COMPONENT MUX_5_TO_1 IS 
		port(
			KEY : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
			X1,X2,X3,X4,X5 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			F : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
		);
	END COMPONENT;
	
	COMPONENT BUFFER_TRI IS 
		port(
			ENTRADA : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
			GATE : IN STD_LOGIC;
			SAIDA: OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
		);
	END COMPONENT;
	
	COMPONENT REG IS 
		port(
			D : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
			R_in,Reset,Clock : IN STD_LOGIC;
			D_out: OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
		);
	END COMPONENT;
	
	COMPONENT REG_BANK IS 
		port(
				REG_READ1,REG_READ2 :IN STD_LOGIC_VECTOR(3 DOWNTO 0);
				WRITE_REG :IN STD_LOGIC_VECTOR(3 DOWNTO 0);
				WRITE_DATA :IN STD_LOGIC_VECTOR(15 DOWNTO 0);
				REG_WRITE: IN STD_LOGIC;
				DATA_READ1 :OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
				DATA_READ2 :OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
				
				R0_OUT : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
				R1_OUT : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
				R2_OUT : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
				R3_OUT : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
				R4_OUT : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
				R5_OUT : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);

				CLOCK : IN STD_LOGIC;
				RESET : IN STD_LOGIC 
		);
	END COMPONENT;
		
	COMPONENT MEMORY is
		 port (
			  ADDRESS  : in  std_logic_vector(15 downto 0);
			  DATA_IN  : in  std_logic_vector(WORD_SIZE-1 downto 0);
			  DATA_OUT : out std_logic_vector(WORD_SIZE-1 downto 0) := (others => '0');
			  READ_MEM : in  std_logic;
			  WRITE_MEM: in  std_logic;
			  CLOCK    : in  std_logic
		 );
	END COMPONENT;
	
			
	COMPONENT INSTRUCTION_MEMORY is
		 port (
			  ADDRESS  : in  std_logic_vector(15 downto 0);
			  DATA_IN  : in  std_logic_vector(WORD_SIZE-1 downto 0);
			  DATA_OUT : out std_logic_vector(WORD_SIZE-1 downto 0) := (others => '0');
			  READ_MEM : in  std_logic;
			  WRITE_MEM: in  std_logic;
			  CLOCK    : in  std_logic
		 );
	END COMPONENT;
	
	COMPONENT TWO_BIT_REG IS 
		port(
			D : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
			R_in,Reset,Clock : IN STD_LOGIC;
			D_out: OUT STD_LOGIC_VECTOR(1 DOWNTO 0)
		);
	END COMPONENT;
	
	COMPONENT SIGN_EXTEND IS 
		 PORT (
			  IN_SIGNAL : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
			  OUT_SIGNAL : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
		 );
	END COMPONENT;
	
	COMPONENT SHIFT_LEFT2 IS 
		PORT (
		  IN_SIGNAL : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		  OUT_SIGNAL : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
		);
	END COMPONENT;
	
	COMPONENT SHIFT_LEFT1 IS 
		PORT (
		  IN_SIGNAL : IN STD_LOGIC_VECTOR(12 DOWNTO 0);
		  OUT_SIGNAL : OUT STD_LOGIC_VECTOR(13 DOWNTO 0)
		);
	END COMPONENT;
	
	COMPONENT PIPE_MEM_WB IS 

	port(
		 -- Inputs
		 MEM_OUT_IN : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 ALU_RESULT_IN : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 IMED_IN : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 REG_DST_IN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);

		 -- Outputs
		 MEM_OUT_OUT : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		 ALU_RESULT_OUT : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		 IMED_OUT : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		 REG_DST_OUT : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);

		 -- Sinais de controle
		 -- WB
		 WB_MEM_TO_REG_IN : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		 WB_REG_WRITE_IN : IN STD_LOGIC;

		 WB_MEM_TO_REG_OUT : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
		 WB_REG_WRITE_OUT : OUT STD_LOGIC;

		 -- Controle de clock e reset
		 CLOCK : IN STD_LOGIC;
		 RESET : IN STD_LOGIC
	);
	END COMPONENT;

	
	COMPONENT PIPE_IF_ID IS 
    port(
        -- Inputs
        NEXT_PC_IN : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
        INSTRUCTION_DATA_IN : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
        IF_ID_WRITE : IN STD_LOGIC;

        -- Outputs
        NEXT_PC_OUT : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
        INSTRUCTION_DATA_OUT : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
        
        -- Sinais de controle de hazard
        IF_FLUSH : IN STD_LOGIC;

        -- Controle de clock e reset
        CLOCK : IN STD_LOGIC;
        RESET : IN STD_LOGIC
    );
	END COMPONENT;
	
COMPONENT PIPE_ID_EX IS 
    port(
        -- Inputs
        A_IN : IN STD_LOGIC_VECTOR(15 DOWNTO 0); -- Registrador A (rs)
        B_IN : IN STD_LOGIC_VECTOR(15 DOWNTO 0); -- Registrador B (rt)
        SIGNAL_EXT_IN : IN STD_LOGIC_VECTOR(15 DOWNTO 0); -- Imediato estendido
        IF_ID_REG_RS_IN : IN STD_LOGIC_VECTOR(3 DOWNTO 0); -- Código do registrador rs
        IF_ID_REG_RT_IN : IN STD_LOGIC_VECTOR(3 DOWNTO 0); -- Código do registrador rt
        IF_ID_REG_RD_IN : IN STD_LOGIC_VECTOR(3 DOWNTO 0); -- Código do registrador rd
        NEXT_PC_IN : IN STD_LOGIC_VECTOR(15 DOWNTO 0); -- Próximo PC

        -- Outputs
        A_OUT : OUT STD_LOGIC_VECTOR(15 DOWNTO 0); -- Registrador A (rs)
        B_OUT : OUT STD_LOGIC_VECTOR(15 DOWNTO 0); -- Registrador B (rt)
        SIGNAL_EXT_OUT : OUT STD_LOGIC_VECTOR(15 DOWNTO 0); -- Imediato estendido
        IF_ID_REG_RS_OUT : OUT STD_LOGIC_VECTOR(3 DOWNTO 0); -- Código do registrador rs
        IF_ID_REG_RT_OUT : OUT STD_LOGIC_VECTOR(3 DOWNTO 0); -- Código do registrador rt
        IF_ID_REG_RD_OUT : OUT STD_LOGIC_VECTOR(3 DOWNTO 0); -- Código do registrador rd
        NEXT_PC_OUT : OUT STD_LOGIC_VECTOR(15 DOWNTO 0); -- Próximo PC

        -- Sinais de controle
        -- EX
        EX_ALU_SRC_IN : IN STD_LOGIC;
        EX_REG_DST_IN : IN STD_LOGIC;
        EX_ALU_OP_IN : IN STD_LOGIC_VECTOR(1 DOWNTO 0);

        EX_ALU_SRC_OUT : OUT STD_LOGIC;
        EX_REG_DST_OUT : OUT STD_LOGIC;
        EX_ALU_OP_OUT : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);

        -- MEM
        MEM_WRITE_IN : IN STD_LOGIC;
        MEM_READ_IN : IN STD_LOGIC;
        -- MEM_ALU_RESULT_IN : IN STD_LOGIC;
        -- MEM_ALU_SRC2_IN : IN STD_LOGIC;

        MEM_WRITE_OUT : OUT STD_LOGIC;
        MEM_READ_OUT : OUT STD_LOGIC;
        -- MEM_ALU_RESULT_OUT : OUT STD_LOGIC;
        -- MEM_ALU_SRC2_OUT : OUT STD_LOGIC;

        -- WB
        WB_MEM_TO_REG_IN : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
        WB_REG_WRITE_IN : IN STD_LOGIC;

        WB_MEM_TO_REG_OUT : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
        WB_REG_WRITE_OUT : OUT STD_LOGIC;

        -- Controle de clock e reset
        CLOCK : IN STD_LOGIC;
        RESET : IN STD_LOGIC

    );
END COMPONENT;

COMPONENT PIPE_EX_MEM IS 

    port(
        -- Inputs
        ALU_OUT_IN : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
        RT_DATA_IN : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
        IMED_IN : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
        REG_DST_IN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);

        -- Outputs
        ALU_OUT_OUT : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);    
        RT_DATA_OUT : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
        IMED_OUT : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
        REG_DST_OUT : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);

        -- Sinais de controle
        -- MEM
        MEM_WRITE_IN : IN STD_LOGIC;
        MEM_READ_IN : IN STD_LOGIC;
        -- MEM_ALU_RESULT_IN : IN STD_LOGIC;
        -- MEM_ALU_SRC2_IN : IN STD_LOGIC;

        MEM_WRITE_OUT : OUT STD_LOGIC;
        MEM_READ_OUT : OUT STD_LOGIC;
        -- MEM_ALU_RESULT_OUT : OUT STD_LOGIC;
        -- MEM_ALU_SRC2_OUT : OUT STD_LOGIC;

        -- WB
        WB_MEM_TO_REG_IN : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
        WB_REG_WRITE_IN : IN STD_LOGIC;

        WB_MEM_TO_REG_OUT : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
        WB_REG_WRITE_OUT : OUT STD_LOGIC;

        -- Controle de clock e reset
        CLOCK : IN STD_LOGIC;
        RESET : IN STD_LOGIC
    );
END COMPONENT;

COMPONENT ONE_BIT_REG IS 
    PORT(
        D      : IN  STD_LOGIC;       -- Entrada de 1 bit
        R_in   : IN  STD_LOGIC;       -- Sinal de controle para escrita
        Reset  : IN  STD_LOGIC;       -- Sinal de reset
        Clock  : IN  STD_LOGIC;       -- Sinal de clock
        D_out  : OUT STD_LOGIC        -- Saída de 1 bit
    );
END COMPONENT;

COMPONENT HAZARD_DETECTION_UNIT IS 
    port(
        PC_WRITE : OUT STD_LOGIC;
        IF_ID_WRITE : OUT STD_LOGIC
    );
END COMPONENT;

COMPONENT FOUR_BIT_REG IS 
	port(
		D : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		R_in,Reset,Clock : IN STD_LOGIC;
		D_out: OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END COMPONENT;


COMPONENT FORWARDING_UNIT IS 
    port(
        RS, RT : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
        
        REG_DST_EX_MEM : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
        REG_DST_MEM_WB : IN STD_LOGIC_VECTOR(3 DOWNTO 0);

        WRITE_REG_EX_MEM : IN STD_LOGIC;
        WRITE_REG_MEM_WB : IN STD_LOGIC;

        FOWARD_A : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
        FOWARD_B : OUT STD_LOGIC_VECTOR(1 DOWNTO 0)
    );
END COMPONENT;

COMPONENT CONTROL_UNIT IS 
    PORT(
        INSTRUCTION : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
        REG_EQUAL : IN STD_LOGIC;

        IF_FLUSH : OUT STD_LOGIC;
        ID_FLUSH : OUT STD_LOGIC;
        EX_FLUSH : OUT STD_LOGIC;
        WB_FLUSH : OUT STD_LOGIC;

        PC_SOURCE : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
        ALU_SRC : OUT STD_LOGIC;
        REG_DST : OUT STD_LOGIC;
        ALU_OP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);

        -- Sinais de controle MEM
        MEM_WRITE : OUT STD_LOGIC;
        MEM_READ : OUT STD_LOGIC;

        -- Sinais de controle WB
        MEM_TO_REG : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
        REG_WRITE : OUT STD_LOGIC;
		  
		  CLOCK : IN STD_LOGIC
    );
END COMPONENT;

COMPONENT ALU_CONTROL IS 
	port(
        ALU_OP  : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
        ADD_SUB : IN STD_LOGIC;
        ALU_CONTROL_OUT : OUT STD_LOGIC
		);
END COMPONENT;
END CPU_PACKAGE;
