LIBRARY ieee;
USE ieee.std_logic_1164.all;
use work.CPU_PACKAGE.all;

ENTITY REG_BANK IS 
	port(
			REG_READ1,REG_READ2 :IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			WRITE_REG :IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			WRITE_DATA :IN STD_LOGIC_VECTOR(15 DOWNTO 0);
			REG_WRITE,REG_READ: IN STD_LOGIC;
			DATA_READ1 :OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
			DATA_READ2 :OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END REG_BANK;

ARCHITECTURE Behavior OF REG_BANK IS
SIGNAL R_IN,WRITE_AUX: STD_LOGIC_VECTOR(0 TO 15);
SIGNAL R0,R1,R2,R3,R4,R5,R6,R7,R8,R9,R10,R11,R12,R13,R14,R15 : STD_LOGIC_VECTOR(3 DOWNTO 0);
BEGIN

	-- Decoder 4 to 16
	WITH WRITE_REG SELECT
		WRITE_AUX <= 	"0000000000000010" WHEN "0001",
						"0000000000000100" WHEN "0010",
						"0000000000001000" WHEN "0011",
						"0000000000010000" WHEN "0100",
						"0000000000100000" WHEN "0101",
						"0000000001000000" WHEN "0110",
						"0000000010000000" WHEN "0111",
						"0000000100000000" WHEN "1000",
						"0000001000000000" WHEN "1001",
						"0000010000000000" WHEN "1010",
						"0000100000000000" WHEN "1011",
						"0001000000000000" WHEN "1100",
						"0010000000000000" WHEN "1101",
						"0100000000000000" WHEN "1110",
						"1000000000000000" WHEN "1111",
						"0000000000000000" WHEN OTHERS;

	
	R_IN(1) <= WRITE_AUX(1) AND REG_WRITE;
	R_IN(2) <= WRITE_AUX(2) AND REG_WRITE;
	R_IN(3) <= WRITE_AUX(3) AND REG_WRITE;
	R_IN(4) <= WRITE_AUX(4) AND REG_WRITE;
	R_IN(5) <= WRITE_AUX(5) AND REG_WRITE;
	R_IN(6) <= WRITE_AUX(6) AND REG_WRITE;
	R_IN(7) <= WRITE_AUX(7) AND REG_WRITE;
	R_IN(8) <= WRITE_AUX(8) AND REG_WRITE;
	R_IN(9) <= WRITE_AUX(9) AND REG_WRITE;
	R_IN(10) <= WRITE_AUX(10) AND REG_WRITE;
	R_IN(11) <= WRITE_AUX(11) AND REG_WRITE;
	R_IN(12) <= WRITE_AUX(12) AND REG_WRITE;
	R_IN(13) <= WRITE_AUX(13) AND REG_WRITE;
	R_IN(14) <= WRITE_AUX(14) AND REG_WRITE;
	R_IN(15) <= WRITE_AUX(15) AND REG_WRITE;

	REG0_INSTANCE: REG PORT MAP("0000000000000000",0,0,CLOCK,R0);
	REG1_INSTANCE: REG PORT MAP(WRITE_DATA,R_in(1),RESET,CLOCK,R1);
	REG2_INSTANCE: REG PORT MAP(WRITE_DATA,R_in(2),RESET,CLOCK,R2);
	REG3_INSTANCE: REG PORT MAP(WRITE_DATA,R_in(3),RESET,CLOCK,R3);
	REG4_INSTANCE: REG PORT MAP(WRITE_DATA,R_in(4),RESET,CLOCK,R4);
	REG5_INSTANCE: REG PORT MAP(WRITE_DATA,R_in(5),RESET,CLOCK,R5);
	REG6_INSTANCE: REG PORT MAP(WRITE_DATA,R_in(6),RESET,CLOCK,R6);
	REG7_INSTANCE: REG PORT MAP(WRITE_DATA,R_in(7),RESET,CLOCK,R7);
	REG8_INSTANCE: REG PORT MAP(WRITE_DATA,R_in(8),RESET,CLOCK,R8);
	REG9_INSTANCE: REG PORT MAP(WRITE_DATA,R_in(9),RESET,CLOCK,R9);
	REG10_INSTANCE: REG PORT MAP(WRITE_DATA,R_in(10),RESET,CLOCK,R10);
	REG11_INSTANCE: REG PORT MAP(WRITE_DATA,R_in(11),RESET,CLOCK,R11);
	REG12_INSTANCE: REG PORT MAP(WRITE_DATA,R_in(12),RESET,CLOCK,R12);
	REG13_INSTANCE: REG PORT MAP(WRITE_DATA,R_in(13),RESET,CLOCK,R13);
	REG14_INSTANCE: REG PORT MAP(WRITE_DATA,R_in(14),RESET,CLOCK,R14);
	REG15_INSTANCE: REG PORT MAP(WRITE_DATA,R_in(15),RESET,CLOCK,R15);

	WITH REG_READ1 SELECT
	MUX1 <= R0 when "0000",
			R1 when "0001",
			R2 when "0010",
			R3 when "0011",
			R4 when "0100",
			R5 when "0101",
			R6 when "0110",
			R7 when "0111",
			R8 when "1000",
			R9 when "1001",
			R10 when "1010",
			R11 when "1011",
			R12 when "1100",
			R13 when "1101",
			R14 when "1110",
			R15 when "1111",
			"0000" when others;

	WITH REG_READ2 SELECT
	MUX2 <= R0 when "0000",
			R1 when "0001",
			R2 when "0010",
			R3 when "0011",
			R4 when "0100",
			R5 when "0101",
			R6 when "0110",
			R7 when "0111",
			R8 when "1000",
			R9 when "1001",
			R10 when "1010",
			R11 when "1011",
			R12 when "1100",
			R13 when "1101",
			R14 when "1110",
			R15 when "1111",
			"0000" when others;
							
	BUFFER1_INSTANCE: BUFFER_TRI PORT MAP(MUX1,REG_READ,DATA_READ1);
	BUFFER2_INSTANCE: BUFFER_TRI PORT MAP(MUX2,REG_READ,DATA_READ2);

END Behavior;
