LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY PIPE_EX_MEM IS 

END PIPE_EX_MEM;
    port(
        ALU_OUT_IN : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
        SECOND_OPERAND_IN : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
        REG_DST_IN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);

        ALU_OUT_OUT : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
        SECOND_OPERAND_OUT : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
        REG_DST_OUT : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
    );

ARCHITECTURE Behavior OF PIPE_EX_MEM IS

BEGIN
END Behavior;
