library ieee;
use ieee.std_logic_1164.all;
USE ieee.STD_LOGIC_unsigned.ALL;

entity UC_LCD is
  port(
	 --Nas entradas ficam todos os sinais que serão observados pela Unidade de controle do display LCD
	 OPCODE : IN STD_LOGIC_VECTOR(7 DOWNTO 0);	
	 CLOCK : IN STD_LOGIC;
	 EQU,GRT,LST,ENABLE : IN STD_LOGIC;
	 
	 -- Nas saídas ficam os sinais de manipulação que controlam o fluxo de dados para o display
	 LCD_DATA : out STD_LOGIC_VECTOR(7 DOWNTO 0); 	-- Palavra de 8-bits para comunicação com o LCD
	 LCD_RW : OUT STD_LOGIC;								-- Sinal para indicar se é leitura ou escrita
	 LCD_EN : OUT STD_LOGIC;								-- Sinal de enable que envia o pulso de comunicação
	 LCD_RS: OUT STD_LOGIC									-- Sinal que indica se é dado ou comando
  );
end entity UC_LCD;

architecture bhv of UC_LCD is

-- Definição de todos os 548 estados da unidade de controle do display LCD
TYPE state_type IS (IDLE_CLEAR1,IDLE_CLEAR2,IDLE,

-- Escrita da primeira linha de cada instrução
SOMA_MSG, SOMA_MSG_EN, SOMA_MSG_TR, SOMA_MENU_MSG, SOMA_MENU_MSG_EN,
SUB_MSG, SUB_MSG_EN, SUB_MSG_TR, SUB_MENU_MSG, SUB_MENU_MSG_EN,
AND_MSG, AND_MSG_EN, AND_MSG_TR, AND_MENU_MSG, AND_MENU_MSG_EN,
OR_MSG, OR_MSG_EN, OR_MSG_TR, OR_MENU_MSG, OR_MENU_MSG_EN,
MUL_MSG, MUL_MSG_EN, MUL_MSG_TR, MUL_MENU_MSG, MUL_MENU_MSG_EN,
NOT_MSG, NOT_MSG_EN, NOT_MSG_TR, NOT_MENU_MSG, NOT_MENU_MSG_EN,
MENU_MSG, MENU_MSG_EN, MENU_MSG_TR,
COMP_MSG, COMP_MSG_EN, COMP_MSG_TR, COMP_MENU_MSG, COMP_MENU_MSG_EN,
LOAD_MSG, LOAD_MSG_EN, LOAD_MSG_TR, LOAD_MENU_MSG, LOAD_MENU_MSG_EN,
SWAP_MSG, SWAP_MSG_EN, SWAP_MSG_TR, SWAP_MENU_MSG, SWAP_MENU_MSG_EN,

-- Estados que gerenciam pooling da segunda linha
SOMA_MENU_X,SOMA_MENU_Y, SOMA_MENU_TRAVA1,SOMA_MENU_TRAVA2,
SUB_MENU_X,SUB_MENU_Y, SUB_MENU_TRAVA1,SUB_MENU_TRAVA2,
AND_MENU_X,AND_MENU_Y, AND_MENU_TRAVA1,AND_MENU_TRAVA2,
OR_MENU_X,OR_MENU_Y, OR_MENU_TRAVA1,OR_MENU_TRAVA2,
MUL_MENU_X,MUL_MENU_Y, MUL_MENU_TRAVA1,MUL_MENU_TRAVA2,
LOAD_MENU_Y, LOAD_MENU_TRAVA1,LOAD_MENU_TRAVA2,
NOT_MENU_X,NOT_MENU_Y, NOT_MENU_TRAVA1,NOT_MENU_TRAVA2,
SWAP_MENU_X,SWAP_MENU_Y, SWAP_MENU_TRAVA1,SWAP_MENU_TRAVA2,
COMP_MENU_X,COMP_MENU_Y,COMP_MENU_OPERATOR, COMP_MENU_TRAVA1,COMP_MENU_TRAVA2,

-- Estados para dar set nos endereços das linhas
LINHA1_ADDRESS_SET,LINHA1_ADDRESS_EN,
LINHA2_ADDRESS_SET,LINHA2_ADDRESS_EN,

-- Escrita da segunda linha da soma
WRITE_RXR1_SOMA,WRITE_RXR1_en_SOMA,WRITE_RXR1_ADDRESS1_SOMA,WRITE_RXR1_1_SOMA,WRITE_RXR1_1_EN_SOMA,WRITE_RXR1_ADDRESS2_SOMA,WRITE_RXR1_ADDRESS2_EN_SOMA,WRITE_1_SOMA,WRITE_1_EN_SOMA,
WRITE_RXR2_SOMA,WRITE_RXR2_en_SOMA,WRITE_RXR2_ADDRESS1_SOMA,WRITE_RXR2_1_SOMA,WRITE_RXR2_1_EN_SOMA,WRITE_RXR2_ADDRESS2_SOMA,WRITE_RXR2_ADDRESS2_EN_SOMA,WRITE_2_SOMA,WRITE_2_EN_SOMA,
WRITE_RXR3_SOMA,WRITE_RXR3_en_SOMA,WRITE_RXR3_ADDRESS1_SOMA,WRITE_RXR3_1_SOMA,WRITE_RXR3_1_EN_SOMA,WRITE_RXR3_ADDRESS2_SOMA,WRITE_RXR3_ADDRESS2_EN_SOMA,WRITE_3_SOMA,WRITE_3_EN_SOMA,
WRITE_RX_SOMA,WRITE_RX_en_SOMA,WRITE_RX_ADDRESS1_SOMA,WRITE_RX_1_SOMA,WRITE_RX_1_EN_SOMA,WRITE_RX_ADDRESS2_SOMA,WRITE_RX_ADDRESS2_EN_SOMA,WRITE_x_SOMA,WRITE_x_EN_SOMA,
WRITE_RYR1_SOMA,WRITE_RYR1_ADDRESS1_SOMA,WRITE_1Y_SOMA,WRITE_1Y_EN_SOMA,
WRITE_RYR2_SOMA,WRITE_RYR2_ADDRESS1_SOMA,WRITE_2Y_SOMA,WRITE_2Y_EN_SOMA,
WRITE_RYR3_SOMA,WRITE_RYR3_ADDRESS1_SOMA,WRITE_3Y_SOMA,WRITE_3Y_EN_SOMA,
WRITE_RY_SOMA,WRITE_RY_ADDRESS1_SOMA,WRITE_Y_SOMA,WRITE_Y_EN_SOMA,

-- Escrita da segunda linha da subtração
WRITE_RXR1_SUB,WRITE_RXR1_en_SUB,WRITE_RXR1_ADDRESS1_SUB,WRITE_RXR1_1_SUB,WRITE_RXR1_1_EN_SUB,WRITE_RXR1_ADDRESS2_SUB,WRITE_RXR1_ADDRESS2_EN_SUB,WRITE_1_SUB,WRITE_1_EN_SUB,
WRITE_RXR2_SUB,WRITE_RXR2_en_SUB,WRITE_RXR2_ADDRESS1_SUB,WRITE_RXR2_1_SUB,WRITE_RXR2_1_EN_SUB,WRITE_RXR2_ADDRESS2_SUB,WRITE_RXR2_ADDRESS2_EN_SUB,WRITE_2_SUB,WRITE_2_EN_SUB,
WRITE_RXR3_SUB,WRITE_RXR3_en_SUB,WRITE_RXR3_ADDRESS1_SUB,WRITE_RXR3_1_SUB,WRITE_RXR3_1_EN_SUB,WRITE_RXR3_ADDRESS2_SUB,WRITE_RXR3_ADDRESS2_EN_SUB,WRITE_3_SUB,WRITE_3_EN_SUB,
WRITE_RX_SUB,WRITE_RX_en_SUB,WRITE_RX_ADDRESS1_SUB,WRITE_RX_1_SUB,WRITE_RX_1_EN_SUB,WRITE_RX_ADDRESS2_SUB,WRITE_RX_ADDRESS2_EN_SUB,WRITE_x_SUB,WRITE_x_EN_SUB,
WRITE_RYR1_SUB,WRITE_RYR1_ADDRESS1_SUB,WRITE_1Y_SUB,WRITE_1Y_EN_SUB,
WRITE_RYR2_SUB,WRITE_RYR2_ADDRESS1_SUB,WRITE_2Y_SUB,WRITE_2Y_EN_SUB,
WRITE_RYR3_SUB,WRITE_RYR3_ADDRESS1_SUB,WRITE_3Y_SUB,WRITE_3Y_EN_SUB,
WRITE_RY_SUB,WRITE_RY_ADDRESS1_SUB,WRITE_Y_SUB,WRITE_Y_EN_SUB,

-- Escrita da segunda linha do AND
WRITE_RXR1_AND,WRITE_RXR1_en_AND,WRITE_RXR1_ADDRESS1_AND,WRITE_RXR1_1_AND,WRITE_RXR1_1_EN_AND,WRITE_RXR1_ADDRESS2_AND,WRITE_RXR1_ADDRESS2_EN_AND,WRITE_1_AND,WRITE_1_EN_AND,
WRITE_RXR2_AND,WRITE_RXR2_en_AND,WRITE_RXR2_ADDRESS1_AND,WRITE_RXR2_1_AND,WRITE_RXR2_1_EN_AND,WRITE_RXR2_ADDRESS2_AND,WRITE_RXR2_ADDRESS2_EN_AND,WRITE_2_AND,WRITE_2_EN_AND,
WRITE_RXR3_AND,WRITE_RXR3_en_AND,WRITE_RXR3_ADDRESS1_AND,WRITE_RXR3_1_AND,WRITE_RXR3_1_EN_AND,WRITE_RXR3_ADDRESS2_AND,WRITE_RXR3_ADDRESS2_EN_AND,WRITE_3_AND,WRITE_3_EN_AND,
WRITE_RX_AND,WRITE_RX_en_AND,WRITE_RX_ADDRESS1_AND,WRITE_RX_1_AND,WRITE_RX_1_EN_AND,WRITE_RX_ADDRESS2_AND,WRITE_RX_ADDRESS2_EN_AND,WRITE_x_AND,WRITE_x_EN_AND,
WRITE_RYR1_AND,WRITE_RYR1_ADDRESS1_AND,WRITE_1Y_AND,WRITE_1Y_EN_AND,
WRITE_RYR2_AND,WRITE_RYR2_ADDRESS1_AND,WRITE_2Y_AND,WRITE_2Y_EN_AND,
WRITE_RYR3_AND,WRITE_RYR3_ADDRESS1_AND,WRITE_3Y_AND,WRITE_3Y_EN_AND,
WRITE_RY_AND,WRITE_RY_ADDRESS1_AND,WRITE_Y_AND,WRITE_Y_EN_AND,

-- Escrita da segunda linha do OR
WRITE_RXR1_OR,WRITE_RXR1_en_OR,WRITE_RXR1_ADDRESS1_OR,WRITE_RXR1_1_OR,WRITE_RXR1_1_EN_OR,WRITE_RXR1_ADDRESS2_OR,WRITE_RXR1_ADDRESS2_EN_OR,WRITE_1_OR,WRITE_1_EN_OR,
WRITE_RXR2_OR,WRITE_RXR2_en_OR,WRITE_RXR2_ADDRESS1_OR,WRITE_RXR2_1_OR,WRITE_RXR2_1_EN_OR,WRITE_RXR2_ADDRESS2_OR,WRITE_RXR2_ADDRESS2_EN_OR,WRITE_2_OR,WRITE_2_EN_OR,
WRITE_RXR3_OR,WRITE_RXR3_en_OR,WRITE_RXR3_ADDRESS1_OR,WRITE_RXR3_1_OR,WRITE_RXR3_1_EN_OR,WRITE_RXR3_ADDRESS2_OR,WRITE_RXR3_ADDRESS2_EN_OR,WRITE_3_OR,WRITE_3_EN_OR,
WRITE_RX_OR,WRITE_RX_en_OR,WRITE_RX_ADDRESS1_OR,WRITE_RX_1_OR,WRITE_RX_1_EN_OR,WRITE_RX_ADDRESS2_OR,WRITE_RX_ADDRESS2_EN_OR,WRITE_x_OR,WRITE_x_EN_OR,
WRITE_RYR1_OR,WRITE_RYR1_ADDRESS1_OR,WRITE_1Y_OR,WRITE_1Y_EN_OR,
WRITE_RYR2_OR,WRITE_RYR2_ADDRESS1_OR,WRITE_2Y_OR,WRITE_2Y_EN_OR,
WRITE_RYR3_OR,WRITE_RYR3_ADDRESS1_OR,WRITE_3Y_OR,WRITE_3Y_EN_OR,
WRITE_RY_OR,WRITE_RY_ADDRESS1_OR,WRITE_Y_OR,WRITE_Y_EN_OR,

-- Escrita da segunda linha da Multiplicação
WRITE_RXR1_MUL,WRITE_RXR1_en_MUL,WRITE_RXR1_ADDRESS1_MUL,WRITE_RXR1_1_MUL,WRITE_RXR1_1_EN_MUL,WRITE_RXR1_ADDRESS2_MUL,WRITE_RXR1_ADDRESS2_EN_MUL,WRITE_1_MUL,WRITE_1_EN_MUL,
WRITE_RXR2_MUL,WRITE_RXR2_en_MUL,WRITE_RXR2_ADDRESS1_MUL,WRITE_RXR2_1_MUL,WRITE_RXR2_1_EN_MUL,WRITE_RXR2_ADDRESS2_MUL,WRITE_RXR2_ADDRESS2_EN_MUL,WRITE_2_MUL,WRITE_2_EN_MUL,
WRITE_RXR3_MUL,WRITE_RXR3_en_MUL,WRITE_RXR3_ADDRESS1_MUL,WRITE_RXR3_1_MUL,WRITE_RXR3_1_EN_MUL,WRITE_RXR3_ADDRESS2_MUL,WRITE_RXR3_ADDRESS2_EN_MUL,WRITE_3_MUL,WRITE_3_EN_MUL,
WRITE_RX_MUL,WRITE_RX_en_MUL,WRITE_RX_ADDRESS1_MUL,WRITE_RX_1_MUL,WRITE_RX_1_EN_MUL,WRITE_RX_ADDRESS2_MUL,WRITE_RX_ADDRESS2_EN_MUL,WRITE_x_MUL,WRITE_x_EN_MUL,
WRITE_RYR1_MUL,WRITE_RYR1_ADDRESS1_MUL,WRITE_1Y_MUL,WRITE_1Y_EN_MUL,
WRITE_RYR2_MUL,WRITE_RYR2_ADDRESS1_MUL,WRITE_2Y_MUL,WRITE_2Y_EN_MUL,
WRITE_RYR3_MUL,WRITE_RYR3_ADDRESS1_MUL,WRITE_3Y_MUL,WRITE_3Y_EN_MUL,
WRITE_RY_MUL,WRITE_RY_ADDRESS1_MUL,WRITE_Y_MUL,WRITE_Y_EN_MUL,

-- Escrita da segunda linha do LOAD
WRITE_RYR1_LOAD,WRITE_RYR1_ADDRESS1_LOAD,WRITE_1Y_LOAD,WRITE_1Y_EN_LOAD,
WRITE_RYR2_LOAD,WRITE_RYR2_ADDRESS1_LOAD,WRITE_2Y_LOAD,WRITE_2Y_EN_LOAD,
WRITE_RYR3_LOAD,WRITE_RYR3_ADDRESS1_LOAD,WRITE_3Y_LOAD,WRITE_3Y_EN_LOAD,
WRITE_RY_LOAD,WRITE_RY_ADDRESS1_LOAD,WRITE_Y_LOAD,WRITE_Y_EN_LOAD,

-- Escrita da segunda linha do NOT
WRITE_RXR1_NOT,WRITE_RXR1_ADDRESS1_NOT,WRITE_RXR1_1_NOT,WRITE_RXR1_1_EN_NOT,
WRITE_RXR2_NOT,WRITE_RXR2_ADDRESS1_NOT,WRITE_RXR2_1_NOT,WRITE_RXR2_1_EN_NOT,
WRITE_RXR3_NOT,WRITE_RXR3_ADDRESS1_NOT,WRITE_RXR3_1_NOT,WRITE_RXR3_1_EN_NOT,
WRITE_RX_NOT,WRITE_RX_ADDRESS1_NOT,WRITE_RX_1_NOT,WRITE_RX_1_EN_NOT,
WRITE_RYR1_NOT,WRITE_RYR1_ADDRESS1_NOT,WRITE_RYR1_1_NOT,WRITE_RYR1_1_EN_NOT,
WRITE_RYR2_NOT,WRITE_RYR2_ADDRESS1_NOT,WRITE_RYR2_1_NOT,WRITE_RYR2_1_EN_NOT,
WRITE_RYR3_NOT,WRITE_RYR3_ADDRESS1_NOT,WRITE_RYR3_1_NOT,WRITE_RYR3_1_EN_NOT,
WRITE_RY_NOT,WRITE_RY_ADDRESS1_NOT,WRITE_RY_1_NOT,WRITE_RY_1_EN_NOT,

-- Escrita da segunda linha do SWAP
WRITE_RXR1_SWAP,WRITE_RXR1_ADDRESS1_SWAP,WRITE_RXR1_1_SWAP,WRITE_RXR1_1_EN_SWAP,
WRITE_RXR2_SWAP,WRITE_RXR2_ADDRESS1_SWAP,WRITE_RXR2_1_SWAP,WRITE_RXR2_1_EN_SWAP,
WRITE_RXR3_SWAP,WRITE_RXR3_ADDRESS1_SWAP,WRITE_RXR3_1_SWAP,WRITE_RXR3_1_EN_SWAP,
WRITE_RX_SWAP,WRITE_RX_ADDRESS1_SWAP,WRITE_RX_1_SWAP,WRITE_RX_1_EN_SWAP,
WRITE_RYR1_SWAP,WRITE_RYR1_ADDRESS1_SWAP,WRITE_RYR1_1_SWAP,WRITE_RYR1_1_EN_SWAP,
WRITE_RYR2_SWAP,WRITE_RYR2_ADDRESS1_SWAP,WRITE_RYR2_1_SWAP,WRITE_RYR2_1_EN_SWAP,
WRITE_RYR3_SWAP,WRITE_RYR3_ADDRESS1_SWAP,WRITE_RYR3_1_SWAP,WRITE_RYR3_1_EN_SWAP,
WRITE_RY_SWAP,WRITE_RY_ADDRESS1_SWAP,WRITE_RY_1_SWAP,WRITE_RY_1_EN_SWAP,

-- Escrita da segunda linha da Comparação
WRITE_RXR1_COMP,WRITE_RXR1_ADDRESS1_COMP,WRITE_RXR1_1_COMP,WRITE_RXR1_1_EN_COMP,
WRITE_RXR2_COMP,WRITE_RXR2_ADDRESS1_COMP,WRITE_RXR2_1_COMP,WRITE_RXR2_1_EN_COMP,
WRITE_RXR3_COMP,WRITE_RXR3_ADDRESS1_COMP,WRITE_RXR3_1_COMP,WRITE_RXR3_1_EN_COMP,
WRITE_RX_COMP,WRITE_RX_ADDRESS1_COMP,WRITE_RX_1_COMP,WRITE_RX_1_EN_COMP,
WRITE_RYR1_COMP,WRITE_RYR1_ADDRESS1_COMP,WRITE_RYR1_1_COMP,WRITE_RYR1_1_EN_COMP,
WRITE_RYR2_COMP,WRITE_RYR2_ADDRESS1_COMP,WRITE_RYR2_1_COMP,WRITE_RYR2_1_EN_COMP,
WRITE_RYR3_COMP,WRITE_RYR3_ADDRESS1_COMP,WRITE_RYR3_1_COMP,WRITE_RYR3_1_EN_COMP,
WRITE_RY_COMP,WRITE_RY_ADDRESS1_COMP,WRITE_RY_1_COMP,WRITE_RY_1_EN_COMP,
COMP_ADDRESS_OPERATOR, COMP_ADDRESS_OPERATOR_EN, COMP_WAIT, COMP_WAIT_EN, COMP_MAIOR, COMP_MAIOR_EN, COMP_MENOR, COMP_MENOR_EN,COMP_IGUAL,COMP_IGUAL_EN

); 
SIGNAL ESTADO : State_type := IDLE_CLEAR1; -- Sinal estado (começa em IDLE_CLEAR1)


SUBTYPE ascii IS STD_LOGIC_VECTOR(7 DOWNTO 0);	-- Este subtipo serve para melhorar a identação dentro dos arrays de mensagens
TYPE CadeiaCaract IS array (1 TO 16) OF ascii;	-- Tipo de array para guardar linha
TYPE init IS ARRAY (1 TO 4) OF ascii;				-- Códigos de iniciação no display

CONSTANT CDG_iniciacao : init:= (x"06",x"0C",x"38",x"01");		-- Códigos de instruções iniciais da placa (CONSULTAR TABELA 6)

-- Vetor para guardar cada linha que será exibida pelo LCD
CONSTANT Linha_SOMA : CadeiaCaract := (x"20",x"20",x"20",x"20",x"20",x"20",x"53",x"4F",x"4D",x"41",x"20",x"20",x"20",x"20",x"20",x"20"); --Inserção de caracteres na primeira linha (array que contém o caractere de cada espaço da primeira linha)
CONSTANT Linha_SUB : CadeiaCaract := (x"20",x"20",x"20",x"53",x"55",x"42",x"54",x"52",x"41",x"43",x"41",x"4F",x"20",x"20",x"20",x"20"); --Inserção de caracteres na primeira linha (array que contém o caractere de cada espaço da primeira linha)
CONSTANT Linha_COMP : CadeiaCaract := (x"20",x"20",x"20",x"43",x"4F",x"4D",x"50",x"41",x"52",x"41",x"43",x"41",x"4F",x"20",x"20",x"20"); --Inserção de caracteres na primeira linha (array que contém o caractere de cada espaço da primeira linha)
CONSTANT Linha_OR : CadeiaCaract := (x"20",x"20",x"20",x"20",x"20",x"41",x"20",x"4F",x"52",x"20",x"42",x"20",x"20",x"20",x"20",x"20"); --Inserção de caracteres na primeira linha (array que contém o caractere de cada espaço da primeira linha)
CONSTANT Linha_AND : CadeiaCaract := (x"20",x"20",x"20",x"20",x"20",x"41",x"20",x"41",x"4E",x"44",x"20",x"42",x"20",x"20",x"20",x"20"); --Inserção de caracteres na primeira linha (array que contém o caractere de cada espaço da primeira linha)
CONSTANT Linha_NOP : CadeiaCaract := (x"20",x"20",x"20",x"20",x"20",x"20",x"4E",x"4F",x"50",x"21",x"20",x"20",x"20",x"20",x"20",x"20"); --Inserção de caracteres na primeira linha (array que contém o caractere de cada espaço da primeira linha)
CONSTANT Linha_MENU : CadeiaCaract := (x"20", x"20", x"20", x"34", x"2D", x"42", x"49", x"54",x"20", x"43", x"50", x"55", x"20", x"20", x"20", x"20");
CONSTANT Linha_NOT : CadeiaCaract := (x"20",x"20",x"20",x"20",x"20",x"4E",x"4F",x"54",x"20",x"42",x"20",x"20",x"20",x"20",x"20",x"20"); --Inserção de caracteres na primeira linha (array que contém o caractere de cada espaço da primeira linha)
CONSTANT Linha_MULT : CadeiaCaract := (x"20", x"4D", x"55", x"4C", x"54", x"49", x"50", x"4C", x"49", x"43", x"41", x"43", x"41", x"4F", x"20", x"20");
CONSTANT Linha_LOAD : CadeiaCaract := (x"20", x"20", x"20", x"20", x"20", x"20", x"4C", x"4F", x"41", x"44", x"20", x"20", x"20", x"20", x"20", x"20");
CONSTANT Linha_SWAP : CadeiaCaract := (x"20", x"20", x"20", x"20", x"20", x"20", x"53", x"57", x"41", x"50", x"20", x"20", x"20", x"20", x"20", x"20");
CONSTANT Linha_MSGOP_SOMA : CadeiaCaract := (x"20", x"20", x"20", x"20", x"52", x"78", x"7F", x"52", x"78", x"2B", x"52", x"79", x"20", x"20", x"20", x"20");
CONSTANT Linha_MSGOP_SUB : CadeiaCaract := (x"20", x"20", x"20", x"20", x"52", x"78", x"7F", x"52", x"78", x"2D", x"52", x"79", x"20", x"20", x"20", x"20");
CONSTANT Linha_MSGOP_MUL : CadeiaCaract := (x"20", x"20", x"20", x"20", x"52", x"78", x"7F", x"52", x"78", x"58", x"52", x"79", x"20", x"20", x"20", x"20");
CONSTANT Linha_MSGOP_AND : CadeiaCaract := (x"20", x"20", x"20", x"20", x"52", x"78", x"7F", x"52", x"78", x"2E", x"52", x"79", x"20", x"20", x"20", x"20");
CONSTANT Linha_MSGOP_OR : CadeiaCaract := (x"20", x"20", x"20", x"20", x"52", x"78", x"7F", x"52", x"78", x"2B", x"52", x"79", x"20", x"20", x"20", x"20");
CONSTANT Linha_MSGOP_LOAD : CadeiaCaract := (x"20", x"20", x"20", x"20", x"52", x"79", x"7F", x"44", x"41", x"54", x"41", x"20", x"20", x"20", x"20", x"20");
CONSTANT Linha_MSGOP_NOT : CadeiaCaract := (x"20", x"20", x"20", x"20", x"20", x"52", x"78", x"7F",x"21", x"52", x"79", x"20", x"20", x"20", x"20", x"20");
CONSTANT Linha_MSGOP_SWAP : CadeiaCaract := (x"20", x"20", x"20", x"20", x"20", x"52", x"78", x"7F", x"7E", x"52", x"79", x"20", x"20", x"20", x"20", x"20");
CONSTANT Linha_MSGOP_COMP : CadeiaCaract := (x"20", x"20", x"20", x"20", x"20", x"52", x"78", x"3F", x"52", x"79", x"20", x"20", x"20", x"20", x"20", x"20");


SIGNAL REG_DATA,OP :STD_LOGIC_VECTOR(3 DOWNTO 0);	-- Sinais auxiliares para melhorar identação
SIGNAL conteiro: INTEGER:=0;								-- Contador que varre as instruções que vâo para o LCD_DATA

BEGIN

-- Instanciando sinais auxiliares
REG_DATA <= OPCODE(3 DOWNTO 0);
OP <= OPCODE(7 DOWNTO 4);

PROCESS (clock)
BEGIN

	IF (clock'EVENT AND clock = '1') THEN
	CASE ESTADO IS
	
		-- ESTADOS IDLE CLEAR RODAM OS COMANDOS DE INICIALIZAÇÃO DO DISPLAY
		WHEN IDLE_CLEAR1 =>
		ESTADO <= IDLE_CLEAR2;
		
		WHEN IDLE_CLEAR2 =>
		conteiro <= conteiro + 1;
		IF conteiro < 4 THEN ESTADO <= IDLE_CLEAR1;
		ELSE ESTADO <= IDLE;
		END IF;
		
		-- ESTADO IDLE É UMA REFERÊNCIA DE "MENU", nele decidimos qual opcde leva a qual mensagem
		WHEN IDLE =>
		conteiro <= 1;
		IF OP = "0000" THEN    ESTADO <= MENU_MSG;--
		ELSIF OP = "0001" THEN ESTADO <= AND_MSG;--
		ELSIF OP = "0010" THEN ESTADO <= OR_MSG;--
		ELSIF OP = "0011" THEN ESTADO <= NOT_MSG;--
		ELSIF OP = "0100" THEN ESTADO <= SOMA_MSG;-- 
		ELSIF OP = "0101" THEN ESTADO <= SUB_MSG;--
		ELSIF OP = "0110" THEN ESTADO <= MUL_MSG;--
		ELSIF OP = "0111" THEN ESTADO <= COMP_MSG;--
		ELSIF OP = "1111" THEN ESTADO <= SWAP_MSG;--
		ELSIF OP = "1000" THEN ESTADO <= LOAD_MSG;--

		ELSE ESTADO <= IDLE;
		END IF;
		
		-- Estado para guiar o cursor para o primeiro caracter da primeira e segunda linha
		WHEN LINHA1_ADDRESS_SET=>
		ESTADO<= LINHA1_ADDRESS_EN;
		
		WHEN LINHA1_ADDRESS_EN=>
		ESTADO <= IDLE;

		
		WHEN LINHA2_ADDRESS_SET=>
		ESTADO<= LINHA2_ADDRESS_EN;
		
		-- Neste estado, precisamos saber qual segunda linha está sendo imprimida
		WHEN LINHA2_ADDRESS_EN=>
		IF OP = "0001" THEN ESTADO <= AND_MENU_MSG;--
		ELSIF OP = "0010" THEN ESTADO <= OR_MENU_MSG;--
		ELSIF OP = "0011" THEN ESTADO <= NOT_MENU_MSG;--
		ELSIF OP = "0100" THEN ESTADO <= SOMA_MENU_MSG;-- 
		ELSIF OP = "0101" THEN ESTADO <= SUB_MENU_MSG;--
		ELSIF OP = "0110" THEN ESTADO <= MUL_MENU_MSG;--
		ELSIF OP = "0111" THEN ESTADO <= COMP_MENU_MSG;--
		ELSIF OP = "1111" THEN ESTADO <= SWAP_MENU_MSG;
		ELSIF OP = "1000" THEN ESTADO <= LOAD_MENU_MSG;--		
		ELSE ESTADO<= LINHA2_ADDRESS_EN;
		END IF;
		
		-- Estados "X_MSG" definem a impressão da primeira linha de cada operação
		WHEN MENU_MSG =>
		ESTADO <= MENU_MSG_EN;
		
		WHEN MENU_MSG_EN =>
		conteiro <= conteiro + 1;
		IF conteiro < 16 THEN ESTADO <= MENU_MSG;
		ELSE ESTADO <= MENU_MSG_TR;
		END IF;
		
		
		WHEN MENU_MSG_TR =>
		conteiro <= 0;
		IF OP = "0000" THEN ESTADO <= MENU_MSG_TR;
		ELSE ESTADO <= LINHA1_ADDRESS_SET;
		END IF;
		
		WHEN LOAD_MSG =>
		ESTADO <= LOAD_MSG_EN;
		
		WHEN LOAD_MSG_EN =>
		conteiro <= conteiro + 1;
		IF conteiro < 16 THEN ESTADO <= LOAD_MSG;
		ELSE ESTADO <= LOAD_MSG_TR;
		END IF;
		
		
		WHEN LOAD_MSG_TR =>
		conteiro <= 1;
		ESTADO <= LINHA2_ADDRESS_SET;

		
		WHEN SWAP_MSG =>
		ESTADO <= SWAP_MSG_EN;
		
		WHEN SWAP_MSG_EN =>
		conteiro <= conteiro + 1;
		IF conteiro < 16 THEN ESTADO <= SWAP_MSG;
		ELSE ESTADO <= SWAP_MSG_TR;
		END IF;
		
		
		WHEN SWAP_MSG_TR =>
		conteiro <= 1;
		ESTADO <= LINHA2_ADDRESS_SET;
		
		WHEN SWAP_MENU_MSG=>
		ESTADO <= SWAP_MENU_MSG_EN;
		
		WHEN SWAP_MENU_MSG_EN=>
		conteiro <= conteiro + 1;
		IF conteiro < 16 THEN ESTADO <= SWAP_MENU_MSG;
		ELSE ESTADO <= SWAP_MENU_X;
		END IF;
		
		
		WHEN SUB_MSG =>
		ESTADO <= SUB_MSG_EN;
		
		WHEN SUB_MSG_EN =>
		conteiro <= conteiro + 1;
		IF conteiro < 16 THEN ESTADO <= SUB_MSG;
		ELSE ESTADO <= SUB_MSG_TR;
		END IF;
		
		
		WHEN SUB_MSG_TR =>
		conteiro <= 1;
		ESTADO <= LINHA2_ADDRESS_SET;
		
		
		WHEN SUB_MENU_MSG=>
		ESTADO <= SUB_MENU_MSG_EN;
		
		WHEN SUB_MENU_MSG_EN=>
		conteiro <= conteiro + 1;
		IF conteiro < 16 THEN ESTADO <= SUB_MENU_MSG;
		ELSE ESTADO <= SUB_MENU_X;
		END IF;
		
		
		
		WHEN MUL_MSG =>
		ESTADO <= MUL_MSG_EN;
		
		WHEN MUL_MSG_EN =>
		conteiro <= conteiro + 1;
		IF conteiro < 16 THEN ESTADO <= MUL_MSG;
		ELSE ESTADO <= MUL_MSG_TR;
		END IF;
		
		
		WHEN MUL_MSG_TR =>
		conteiro <= 1;
		ESTADO <= LINHA2_ADDRESS_SET;
		
		
		WHEN MUL_MENU_MSG=>
		ESTADO <= MUL_MENU_MSG_EN;
		
		WHEN MUL_MENU_MSG_EN=>
		conteiro <= conteiro + 1;
		IF conteiro < 16 THEN ESTADO <= MUL_MENU_MSG;
		ELSE ESTADO <= MUL_MENU_X;
		END IF;
		
		
		
		WHEN AND_MSG =>
		ESTADO <= AND_MSG_EN;
		
		WHEN AND_MSG_EN =>
		conteiro <= conteiro + 1;
		IF conteiro < 16 THEN ESTADO <= AND_MSG;
		ELSE ESTADO <= AND_MSG_TR;
		END IF;
		
		
		WHEN AND_MSG_TR =>
		conteiro <= 1;
		ESTADO <= LINHA2_ADDRESS_SET;
		
		
		WHEN AND_MENU_MSG=>
		ESTADO <= AND_MENU_MSG_EN;
		
		WHEN AND_MENU_MSG_EN=>
		conteiro <= conteiro + 1;
		IF conteiro < 16 THEN ESTADO <= AND_MENU_MSG;
		ELSE ESTADO <= AND_MENU_X;
		END IF;
		
		
		
		WHEN OR_MSG =>
		ESTADO <= OR_MSG_EN;
		
		WHEN OR_MSG_EN =>
		conteiro <= conteiro + 1;
		IF conteiro < 16 THEN ESTADO <= OR_MSG;
		ELSE ESTADO <= OR_MSG_TR;
		END IF;
		
		
		WHEN OR_MSG_TR =>
		conteiro <= 1;
		ESTADO <= LINHA2_ADDRESS_SET;
		
		
		WHEN OR_MENU_MSG=>
		ESTADO <= OR_MENU_MSG_EN;
		
		WHEN OR_MENU_MSG_EN=>
		conteiro <= conteiro + 1;
		IF conteiro < 16 THEN ESTADO <= OR_MENU_MSG;
		ELSE ESTADO <= OR_MENU_X;
		END IF;
		
		
		
		WHEN NOT_MSG =>
		ESTADO <= NOT_MSG_EN;
		
		WHEN NOT_MSG_EN =>
		conteiro <= conteiro + 1;
		IF conteiro < 16 THEN ESTADO <= NOT_MSG;
		ELSE ESTADO <= NOT_MSG_TR;
		END IF;
		
		
		WHEN NOT_MSG_TR =>
		conteiro <= 1;
		ESTADO <= LINHA2_ADDRESS_SET;
		
		WHEN NOT_MENU_MSG=>
		ESTADO <= NOT_MENU_MSG_EN;
		
		WHEN NOT_MENU_MSG_EN=>
		conteiro <= conteiro + 1;
		IF conteiro < 16 THEN ESTADO <= NOT_MENU_MSG;
		ELSE ESTADO <= NOT_MENU_X;
		END IF;
		
		WHEN COMP_MSG =>
		ESTADO <= COMP_MSG_EN;
		
		WHEN COMP_MSG_EN =>
		conteiro <= conteiro + 1;
		IF conteiro < 16 THEN ESTADO <= COMP_MSG;
		ELSE ESTADO <= COMP_MSG_TR;
		END IF;
		
		
		WHEN COMP_MSG_TR =>
		conteiro <= 1;
		ESTADO <= LINHA2_ADDRESS_SET;
		
		WHEN COMP_MENU_MSG=>
		ESTADO <= COMP_MENU_MSG_EN;
		
		WHEN COMP_MENU_MSG_EN=>
		conteiro <= conteiro + 1;
		IF conteiro < 16 THEN ESTADO <= COMP_MENU_MSG;
		ELSE ESTADO <= COMP_MENU_X;
		END IF;
		
----------------------------------------------------------

		WHEN SOMA_MSG =>
		ESTADO <= SOMA_MSG_EN;
		
		WHEN SOMA_MSG_EN =>
		conteiro <= conteiro + 1;
		IF conteiro < 16 THEN ESTADO <= SOMA_MSG;
		ELSE ESTADO <= SOMA_MSG_TR;
		END IF;
		
		
		WHEN SOMA_MSG_TR =>
		conteiro <= 1;
		ESTADO <= LINHA2_ADDRESS_SET;
		
		
		WHEN SOMA_MENU_MSG=>
		ESTADO <= SOMA_MENU_MSG_EN;
		
		WHEN SOMA_MENU_MSG_EN=>
		conteiro <= conteiro + 1;
		IF conteiro < 16 THEN ESTADO <= SOMA_MENU_MSG;
		ELSE ESTADO <= SOMA_MENU_X;
		END IF;
		
		-- Estados "X_MENU_X" indicam o estado que faz a interpretação da segunda parte do OPCODE,
		-- nele decidimos se vamos imprimir "1,2,3,x ou y" na segunda parte da mensagem
		WHEN SOMA_MENU_X=>
		conteiro <= 0;
		
		IF (REG_DATA(3 DOWNTO 2) = "01") AND (OP="0100") THEN
		ESTADO <= WRITE_RXR1_SOMA;
		
		ELSIF REG_DATA(3 DOWNTO 2) = "10" AND (OP="0100")THEN
		ESTADO <= WRITE_RXR2_SOMA;
--		
		ELSIF REG_DATA(3 DOWNTO 2) = "11" AND (OP="0100")THEN
		ESTADO <= WRITE_RXR3_SOMA;
		
		ELSIF REG_DATA(3 DOWNTO 2) = "00" AND (OP="0100")THEN
		ESTADO <= WRITE_RX_SOMA;
		
		ELSE
		ESTADO <=SOMA_MENU_TRAVA1;
		END IF;
				
				
				
		WHEN SOMA_MENU_Y=>
		IF REG_DATA(1 DOWNTO 0) = "01" AND (OP="0100")THEN
		ESTADO <= WRITE_RYR1_SOMA;
		
		ELSIF REG_DATA(1 DOWNTO 0) = "10" AND (OP="0100")THEN
		ESTADO <= WRITE_RYR2_SOMA;
		
		ELSIF REG_DATA(1 DOWNTO 0) = "11" AND (OP="0100") THEN
		ESTADO <= WRITE_RYR3_SOMA;
		
		ELSIF REG_DATA(1 DOWNTO 0) = "00" AND (OP="0100")THEN
		ESTADO <= WRITE_RY_SOMA;
		
		ELSE
		ESTADO <=SOMA_MENU_TRAVA1;
		
		END IF;
		
		
		WHEN SOMA_MENU_TRAVA1 =>
		IF OP="0100" THEN
		ESTADO <= SOMA_MENU_X;
		ELSE 	ESTADO <= SOMA_MENU_TRAVA2;
		END IF;

		WHEN SOMA_MENU_TRAVA2 =>
		IF NOT OP="0100" THEN
		ESTADO <= SOMA_MENU_X;
		ELSE 	ESTADO <= IDLE_CLEAR1;
		END IF;
		
		
		
		
		WHEN SUB_MENU_X=>
		conteiro <= 0;
		
		IF (REG_DATA(3 DOWNTO 2) = "01") AND (OP="0101") THEN
		ESTADO <= WRITE_RXR1_SUB;
		
		ELSIF REG_DATA(3 DOWNTO 2) = "10" AND (OP="0101")THEN
		ESTADO <= WRITE_RXR2_SUB;
--		
		ELSIF REG_DATA(3 DOWNTO 2) = "11" AND (OP="0101")THEN
		ESTADO <= WRITE_RXR3_SUB;
		
		ELSIF REG_DATA(3 DOWNTO 2) = "00" AND (OP="0101")THEN
		ESTADO <= WRITE_RX_SUB;
		
		ELSE
		ESTADO <=SUB_MENU_TRAVA1;
		END IF;
				
				
				
		WHEN SUB_MENU_Y=>
		IF REG_DATA(1 DOWNTO 0) = "01" AND (OP="0101")THEN
		ESTADO <= WRITE_RYR1_SUB;
		
		ELSIF REG_DATA(1 DOWNTO 0) = "10" AND (OP="0101")THEN
		ESTADO <= WRITE_RYR2_SUB;
		
		ELSIF REG_DATA(1 DOWNTO 0) = "11" AND (OP="0101") THEN
		ESTADO <= WRITE_RYR3_SUB;
		
		ELSIF REG_DATA(1 DOWNTO 0) = "00" AND (OP="0101")THEN
		ESTADO <= WRITE_RY_SUB;
		
		ELSE
		ESTADO <=SUB_MENU_TRAVA1;
		
		END IF;
		
		
		WHEN SUB_MENU_TRAVA1 =>
		IF OP="0101" THEN
		ESTADO <= SUB_MENU_X;
		ELSE 	ESTADO <= SUB_MENU_TRAVA2;
		END IF;

		WHEN SUB_MENU_TRAVA2 =>
		IF NOT OP="0101" THEN
		ESTADO <= SUB_MENU_X;
		ELSE 	ESTADO <= IDLE_CLEAR1;
		END IF;
		
		
		WHEN AND_MENU_X=>
		conteiro <= 0;
		
		IF (REG_DATA(3 DOWNTO 2) = "01") AND (OP="0001") THEN
		ESTADO <= WRITE_RXR1_AND;
		
		ELSIF REG_DATA(3 DOWNTO 2) = "10" AND (OP="0001")THEN
		ESTADO <= WRITE_RXR2_AND;
--		
		ELSIF REG_DATA(3 DOWNTO 2) = "11" AND (OP="0001")THEN
		ESTADO <= WRITE_RXR3_AND;
		
		ELSIF REG_DATA(3 DOWNTO 2) = "00" AND (OP="0001")THEN
		ESTADO <= WRITE_RX_AND;
		
		ELSE
		ESTADO <=AND_MENU_TRAVA1;
		END IF;
				
				
				
		WHEN AND_MENU_Y=>
		IF REG_DATA(1 DOWNTO 0) = "01" AND (OP="0001")THEN
		ESTADO <= WRITE_RYR1_AND;
		
		ELSIF REG_DATA(1 DOWNTO 0) = "10" AND (OP="0001")THEN
		ESTADO <= WRITE_RYR2_AND;
		
		ELSIF REG_DATA(1 DOWNTO 0) = "11" AND (OP="0001") THEN
		ESTADO <= WRITE_RYR3_AND;
		
		ELSIF REG_DATA(1 DOWNTO 0) = "00" AND (OP="0001")THEN
		ESTADO <= WRITE_RY_AND;
		
		ELSE
		ESTADO <=AND_MENU_TRAVA1;
		
		END IF;
		
		
		WHEN AND_MENU_TRAVA1 =>
		IF OP="0101" THEN
		ESTADO <= AND_MENU_X;
		ELSE 	ESTADO <= AND_MENU_TRAVA2;
		END IF;

		WHEN AND_MENU_TRAVA2 =>
		IF NOT OP="0101" THEN
		ESTADO <= AND_MENU_X;
		ELSE 	ESTADO <= IDLE_CLEAR1;
		END IF;
	
	
	
		WHEN OR_MENU_X=>
		conteiro <= 0;
		
		IF (REG_DATA(3 DOWNTO 2) = "01") AND (OP="0010") THEN
		ESTADO <= WRITE_RXR1_OR;
		
		ELSIF REG_DATA(3 DOWNTO 2) = "10" AND (OP="0010")THEN
		ESTADO <= WRITE_RXR2_OR;
--		
		ELSIF REG_DATA(3 DOWNTO 2) = "11" AND (OP="0010")THEN
		ESTADO <= WRITE_RXR3_OR;
		
		ELSIF REG_DATA(3 DOWNTO 2) = "00" AND (OP="0010")THEN
		ESTADO <= WRITE_RX_OR;
		
		ELSE
		ESTADO <=OR_MENU_TRAVA1;
		END IF;
				
				
				
		WHEN OR_MENU_Y=>
		IF REG_DATA(1 DOWNTO 0) = "01" AND (OP="0010")THEN
		ESTADO <= WRITE_RYR1_OR;
		
		ELSIF REG_DATA(1 DOWNTO 0) = "10" AND (OP="0010")THEN
		ESTADO <= WRITE_RYR2_OR;
		
		ELSIF REG_DATA(1 DOWNTO 0) = "11" AND (OP="0010") THEN
		ESTADO <= WRITE_RYR3_OR;
		
		ELSIF REG_DATA(1 DOWNTO 0) = "00" AND (OP="0010")THEN
		ESTADO <= WRITE_RY_OR;
		
		ELSE
		ESTADO <=OR_MENU_TRAVA1;
		
		END IF;
		
		
		WHEN OR_MENU_TRAVA1 =>
		IF OP="0010" THEN
		ESTADO <= OR_MENU_X;
		ELSE 	ESTADO <= OR_MENU_TRAVA2;
		END IF;

		WHEN OR_MENU_TRAVA2 =>
		IF NOT OP="0010" THEN
		ESTADO <= OR_MENU_X;
		ELSE 	ESTADO <= IDLE_CLEAR1;
		END IF;
		
		
		WHEN MUL_MENU_X=>
		conteiro <= 0;
		
		IF (REG_DATA(3 DOWNTO 2) = "01") AND (OP="0110") THEN
		ESTADO <= WRITE_RXR1_MUL;
		
		ELSIF REG_DATA(3 DOWNTO 2) = "10" AND (OP="0110")THEN
		ESTADO <= WRITE_RXR2_MUL;
--		
		ELSIF REG_DATA(3 DOWNTO 2) = "11" AND (OP="0110")THEN
		ESTADO <= WRITE_RXR3_MUL;
		
		ELSIF REG_DATA(3 DOWNTO 2) = "00" AND (OP="0110")THEN
		ESTADO <= WRITE_RX_MUL;
		
		ELSE
		ESTADO <=MUL_MENU_TRAVA1;
		END IF;
				
				
				
		WHEN MUL_MENU_Y=>
		IF REG_DATA(1 DOWNTO 0) = "01" AND (OP="0110")THEN
		ESTADO <= WRITE_RYR1_MUL;
		
		ELSIF REG_DATA(1 DOWNTO 0) = "10" AND (OP="0110")THEN
		ESTADO <= WRITE_RYR2_MUL;
		
		ELSIF REG_DATA(1 DOWNTO 0) = "11" AND (OP="0110") THEN
		ESTADO <= WRITE_RYR3_MUL;
		
		ELSIF REG_DATA(1 DOWNTO 0) = "00" AND (OP="0110")THEN
		ESTADO <= WRITE_RY_MUL;
		
		ELSE
		ESTADO <=MUL_MENU_TRAVA1;
		
		END IF;
		
		
		WHEN MUL_MENU_TRAVA1 =>
		IF OP="0110" THEN
		ESTADO <= MUL_MENU_X;
		ELSE 	ESTADO <= MUL_MENU_TRAVA2;
		END IF;

		WHEN MUL_MENU_TRAVA2 =>
		IF NOT OP="0110" THEN
		ESTADO <= MUL_MENU_X;
		ELSE 	ESTADO <= IDLE_CLEAR1;
		END IF;


		WHEN LOAD_MENU_MSG=>
		ESTADO <= LOAD_MENU_MSG_EN;
		
		WHEN LOAD_MENU_MSG_EN=>
		conteiro <= conteiro + 1;
		IF conteiro < 16 THEN ESTADO <= LOAD_MENU_MSG;
		ELSE ESTADO <= LOAD_MENU_Y;
		END IF;
		
		WHEN LOAD_MENU_Y=>
		conteiro <= 0;
		
		IF (REG_DATA(1 DOWNTO 0) = "01") AND (OP="1000") THEN
		ESTADO <= WRITE_RYR1_LOAD;
		
		ELSIF REG_DATA(1 DOWNTO 0) = "10" AND (OP="1000")THEN
		ESTADO <= WRITE_RYR2_LOAD;
--		
		ELSIF REG_DATA(1 DOWNTO 0) = "11" AND (OP="1000")THEN
		ESTADO <= WRITE_RYR3_LOAD;
		
		ELSIF REG_DATA(1 DOWNTO 0) = "00" AND (OP="1000")THEN
		ESTADO <= WRITE_RY_LOAD;
		
		ELSE
		ESTADO <=LOAD_MENU_TRAVA1;
		END IF;
				
		
		
		WHEN LOAD_MENU_TRAVA1 =>
		IF OP="1000" THEN
		ESTADO <= LOAD_MENU_Y;
		ELSE 	ESTADO <= LOAD_MENU_TRAVA2;
		END IF;

		WHEN LOAD_MENU_TRAVA2 =>
		IF NOT OP="1000" THEN
		ESTADO <= LOAD_MENU_Y;
		ELSE 	ESTADO <= IDLE_CLEAR1;
		END IF;
		
		
		WHEN NOT_MENU_X=>
		conteiro <= 0;
		
		IF (REG_DATA(3 DOWNTO 2) = "01") AND (OP="0011") THEN
		ESTADO <= WRITE_RXR1_NOT;
		
		ELSIF REG_DATA(3 DOWNTO 2) = "10" AND (OP="0011")THEN
		ESTADO <= WRITE_RXR2_NOT;
--		
		ELSIF REG_DATA(3 DOWNTO 2) = "11" AND (OP="0011")THEN
		ESTADO <= WRITE_RXR3_NOT;
		
		ELSIF REG_DATA(3 DOWNTO 2) = "00" AND (OP="0011")THEN
		ESTADO <= WRITE_RX_NOT;
		
		ELSE
		ESTADO <=NOT_MENU_TRAVA1;
		END IF;
				
				
				
		WHEN NOT_MENU_Y=>
		IF REG_DATA(1 DOWNTO 0) = "01" AND (OP="0011")THEN
		ESTADO <= WRITE_RYR1_NOT;
		
		ELSIF REG_DATA(1 DOWNTO 0) = "10" AND (OP="0011")THEN
		ESTADO <= WRITE_RYR2_NOT;
		
		ELSIF REG_DATA(1 DOWNTO 0) = "11" AND (OP="0011") THEN
		ESTADO <= WRITE_RYR3_NOT;
		
		ELSIF REG_DATA(1 DOWNTO 0) = "00" AND (OP="0011")THEN
		ESTADO <= WRITE_RY_NOT;
		
		ELSE
		ESTADO <=NOT_MENU_TRAVA1;
		
		END IF;
		
		
		WHEN NOT_MENU_TRAVA1 =>
		IF OP="0011" THEN
		ESTADO <= NOT_MENU_X;
		ELSE 	ESTADO <= NOT_MENU_TRAVA2;
		END IF;

		WHEN NOT_MENU_TRAVA2 =>
		IF NOT OP="0011" THEN
		ESTADO <= NOT_MENU_X;
		ELSE 	ESTADO <= IDLE_CLEAR1;
		END IF;
		
		
		
		
		WHEN SWAP_MENU_X=>
		conteiro <= 0;
		
		IF (REG_DATA(3 DOWNTO 2) = "01") AND (OP="1111") THEN
		ESTADO <= WRITE_RXR1_SWAP;
		
		ELSIF REG_DATA(3 DOWNTO 2) = "10" AND (OP="1111")THEN
		ESTADO <= WRITE_RXR2_SWAP;
--		
		ELSIF REG_DATA(3 DOWNTO 2) = "11" AND (OP="1111")THEN
		ESTADO <= WRITE_RXR3_SWAP;
		
		ELSIF REG_DATA(3 DOWNTO 2) = "00" AND (OP="1111")THEN
		ESTADO <= WRITE_RX_SWAP;
		
		ELSE
		ESTADO <=SWAP_MENU_TRAVA1;
		END IF;
				
				
				
		WHEN SWAP_MENU_Y=>
		IF REG_DATA(1 DOWNTO 0) = "01" AND (OP="1111")THEN
		ESTADO <= WRITE_RYR1_SWAP;
		
		ELSIF REG_DATA(1 DOWNTO 0) = "10" AND (OP="1111")THEN
		ESTADO <= WRITE_RYR2_SWAP;
		
		ELSIF REG_DATA(1 DOWNTO 0) = "11" AND (OP="1111") THEN
		ESTADO <= WRITE_RYR3_SWAP;
		
		ELSIF REG_DATA(1 DOWNTO 0) = "00" AND (OP="1111")THEN
		ESTADO <= WRITE_RY_SWAP;
		
		ELSE
		ESTADO <=SWAP_MENU_TRAVA1;
		
		END IF;
		
		
		WHEN SWAP_MENU_TRAVA1 =>
		IF OP="1111" THEN
		ESTADO <= SWAP_MENU_X;
		ELSE 	ESTADO <= SWAP_MENU_TRAVA2;
		END IF;

		WHEN SWAP_MENU_TRAVA2 =>
		IF NOT OP="1111" THEN
		ESTADO <= SWAP_MENU_X;
		ELSE 	ESTADO <= IDLE_CLEAR1;
		END IF;
		
		
		WHEN COMP_MENU_X=>
		conteiro <= 0;
		
		IF (REG_DATA(3 DOWNTO 2) = "01") AND (OP="0111") THEN
		ESTADO <= WRITE_RXR1_COMP;
		
		ELSIF REG_DATA(3 DOWNTO 2) = "10" AND (OP="0111")THEN
		ESTADO <= WRITE_RXR2_COMP;
--		
		ELSIF REG_DATA(3 DOWNTO 2) = "11" AND (OP="0111")THEN
		ESTADO <= WRITE_RXR3_COMP;
		
		ELSIF REG_DATA(3 DOWNTO 2) = "00" AND (OP="0111")THEN
		ESTADO <= WRITE_RX_COMP;
		
		ELSE
		ESTADO <=COMP_MENU_TRAVA1;
		END IF;
				
				
				
		WHEN COMP_MENU_Y=>
		IF REG_DATA(1 DOWNTO 0) = "01" AND (OP="0111")THEN
		ESTADO <= WRITE_RYR1_COMP;
		
		ELSIF REG_DATA(1 DOWNTO 0) = "10" AND (OP="0111")THEN
		ESTADO <= WRITE_RYR2_COMP;
		
		ELSIF REG_DATA(1 DOWNTO 0) = "11" AND (OP="0111") THEN
		ESTADO <= WRITE_RYR3_COMP;
		
		ELSIF REG_DATA(1 DOWNTO 0) = "00" AND (OP="0111")THEN
		ESTADO <= WRITE_RY_COMP;
		
		ELSE
		ESTADO <=COMP_MENU_TRAVA1;
		
		END IF;
		
		WHEN COMP_MENU_OPERATOR =>
		ESTADO <= COMP_ADDRESS_OPERATOR;
		
		WHEN COMP_MENU_TRAVA1 =>
		IF OP="0111" THEN
		ESTADO <= COMP_MENU_X;
		ELSE 	ESTADO <= COMP_MENU_TRAVA2;
		END IF;

		WHEN COMP_MENU_TRAVA2 =>
		IF NOT OP="0111" THEN
		ESTADO <= COMP_MENU_X;
		ELSE 	ESTADO <= IDLE_CLEAR1;
		END IF;		
		

-----------------------------------------------------------------

-- Essas sequencias de estados servem para alinhar os endereços dos caracteres solicitados no
-- estado anterior com seus respectivos endereços para todos os casos em todas as intruçoes

		WHEN WRITE_RXR1_SOMA=>
		ESTADO<=WRITE_RXR1_ADDRESS1_SOMA;
		
		WHEN WRITE_RXR1_ADDRESS1_SOMA=>
		ESTADO<= WRITE_RXR1_1_SOMA;
		
		WHEN WRITE_RXR1_1_SOMA=>
		ESTADO<= WRITE_RXR1_1_EN_SOMA;
		
		WHEN WRITE_RXR1_1_EN_SOMA=>
		ESTADO<= WRITE_RXR1_ADDRESS2_SOMA;
		
		WHEN WRITE_RXR1_ADDRESS2_SOMA=>
		ESTADO<= WRITE_RXR1_ADDRESS2_EN_SOMA;
		
		WHEN WRITE_RXR1_ADDRESS2_EN_SOMA=>
		ESTADO<= WRITE_1_SOMA;
		
		WHEN WRITE_1_SOMA=>
		ESTADO <= WRITE_1_EN_SOMA;
		
		WHEN WRITE_1_EN_SOMA =>
		ESTADO<= SOMA_MENU_Y;

		
		WHEN WRITE_RXR2_SOMA=>
		ESTADO<=WRITE_RXR2_ADDRESS1_SOMA;
		
		WHEN WRITE_RXR2_ADDRESS1_SOMA=>
		ESTADO<= WRITE_RXR2_1_SOMA;
		
		WHEN WRITE_RXR2_1_SOMA=>
		ESTADO<= WRITE_RXR2_1_EN_SOMA;
		
		WHEN WRITE_RXR2_1_EN_SOMA=>
		ESTADO<= WRITE_RXR2_ADDRESS2_SOMA;
		
		WHEN WRITE_RXR2_ADDRESS2_SOMA=>
		ESTADO<= WRITE_RXR2_ADDRESS2_EN_SOMA;
		
		WHEN WRITE_RXR2_ADDRESS2_EN_SOMA=>
		ESTADO<= WRITE_2_SOMA;
		
		WHEN WRITE_2_SOMA=>
		ESTADO <= WRITE_2_EN_SOMA;
		
		WHEN WRITE_2_EN_SOMA =>	
		ESTADO<= SOMA_MENU_Y;
	
		
		WHEN WRITE_RXR3_SOMA=>
		ESTADO<=WRITE_RXR3_ADDRESS1_SOMA;
		
		WHEN WRITE_RXR3_ADDRESS1_SOMA=>
		ESTADO<= WRITE_RXR3_1_SOMA;
		
		WHEN WRITE_RXR3_1_SOMA=>
		ESTADO<= WRITE_RXR3_1_EN_SOMA;
		
		WHEN WRITE_RXR3_1_EN_SOMA=>
		ESTADO<= WRITE_RXR3_ADDRESS2_SOMA;
		
		WHEN WRITE_RXR3_ADDRESS2_SOMA=>
		ESTADO<= WRITE_RXR3_ADDRESS2_EN_SOMA;
		
		WHEN WRITE_RXR3_ADDRESS2_EN_SOMA=>
		ESTADO<= WRITE_3_SOMA;
		
		WHEN WRITE_3_SOMA=>
		ESTADO <= WRITE_3_EN_SOMA;
		
		WHEN WRITE_3_EN_SOMA =>
		ESTADO<= SOMA_MENU_Y;
	
		
		WHEN WRITE_RX_SOMA=>
		ESTADO<=WRITE_RX_ADDRESS1_SOMA;
		
		WHEN WRITE_RX_ADDRESS1_SOMA=>
		ESTADO<= WRITE_RX_1_SOMA;
		
		WHEN WRITE_RX_1_SOMA=>
		ESTADO<= WRITE_RX_1_EN_SOMA;
		
		WHEN WRITE_RX_1_EN_SOMA=>
		ESTADO<= WRITE_RX_ADDRESS2_SOMA;
		
		WHEN WRITE_RX_ADDRESS2_SOMA=>
		ESTADO<= WRITE_RX_ADDRESS2_EN_SOMA;
		
		WHEN WRITE_RX_ADDRESS2_EN_SOMA=>
		ESTADO<= WRITE_x_SOMA;
		
		WHEN WRITE_x_SOMA=>
		ESTADO <= WRITE_x_EN_SOMA;
		
		WHEN WRITE_x_EN_SOMA =>	
		ESTADO<= SOMA_MENU_Y;
		
		
		
		

		WHEN WRITE_RYR1_SOMA=>
		ESTADO<=WRITE_RYR1_ADDRESS1_SOMA;
		
		WHEN WRITE_RYR1_ADDRESS1_SOMA=>
		ESTADO<= WRITE_1Y_SOMA;
		
		WHEN WRITE_1Y_SOMA=>
		ESTADO <= WRITE_1Y_EN_SOMA;
		
		WHEN WRITE_1Y_EN_SOMA =>
		ESTADO<= SOMA_MENU_X;

		
		WHEN WRITE_RYR2_SOMA=>
		ESTADO<=WRITE_RYR2_ADDRESS1_SOMA;
		
		WHEN WRITE_RYR2_ADDRESS1_SOMA=>
		ESTADO<= WRITE_2Y_SOMA;
		
		WHEN WRITE_2Y_SOMA=>
		ESTADO <= WRITE_2Y_EN_SOMA;
		
		WHEN WRITE_2Y_EN_SOMA =>
		ESTADO<= SOMA_MENU_X;
	
	
		
		WHEN WRITE_RYR3_SOMA=>
		ESTADO<=WRITE_RYR3_ADDRESS1_SOMA;
		
		WHEN WRITE_RYR3_ADDRESS1_SOMA=>
		ESTADO<= WRITE_3Y_SOMA;
		
		WHEN WRITE_3Y_SOMA=>
		ESTADO <= WRITE_3Y_EN_SOMA;
		
		WHEN WRITE_3Y_EN_SOMA =>
		ESTADO<= SOMA_MENU_X;
			
		
		WHEN WRITE_RY_SOMA=>
		ESTADO<=WRITE_RY_ADDRESS1_SOMA;
		
		WHEN WRITE_RY_ADDRESS1_SOMA=>
		ESTADO<= WRITE_Y_SOMA;
		
		WHEN WRITE_Y_SOMA=>
		ESTADO <= WRITE_Y_EN_SOMA;
		
		WHEN WRITE_Y_EN_SOMA =>
		ESTADO<= SOMA_MENU_X;
		

---------------------------------------------------------------
---------------------------------------------------------------
		
		
		WHEN WRITE_RXR1_SUB=>
		ESTADO<=WRITE_RXR1_ADDRESS1_SUB;
		
		WHEN WRITE_RXR1_ADDRESS1_SUB=>
		ESTADO<= WRITE_RXR1_1_SUB;
		
		WHEN WRITE_RXR1_1_SUB=>
		ESTADO<= WRITE_RXR1_1_EN_SUB;
		
		WHEN WRITE_RXR1_1_EN_SUB=>
		ESTADO<= WRITE_RXR1_ADDRESS2_SUB;
		
		WHEN WRITE_RXR1_ADDRESS2_SUB=>
		ESTADO<= WRITE_RXR1_ADDRESS2_EN_SUB;
		
		WHEN WRITE_RXR1_ADDRESS2_EN_SUB=>
		ESTADO<= WRITE_1_SUB;
		
		WHEN WRITE_1_SUB=>
		ESTADO <= WRITE_1_EN_SUB;
		
		WHEN WRITE_1_EN_SUB =>
		ESTADO<= SUB_MENU_Y;
		
		
		WHEN WRITE_RXR2_SUB=>
		ESTADO<=WRITE_RXR2_ADDRESS1_SUB;
		
		WHEN WRITE_RXR2_ADDRESS1_SUB=>
		ESTADO<= WRITE_RXR2_1_SUB;
		
		WHEN WRITE_RXR2_1_SUB=>
		ESTADO<= WRITE_RXR2_1_EN_SUB;
		
		WHEN WRITE_RXR2_1_EN_SUB=>
		ESTADO<= WRITE_RXR2_ADDRESS2_SUB;
		
		WHEN WRITE_RXR2_ADDRESS2_SUB=>
		ESTADO<= WRITE_RXR2_ADDRESS2_EN_SUB;
		
		WHEN WRITE_RXR2_ADDRESS2_EN_SUB=>
		ESTADO<= WRITE_2_SUB;
		
		WHEN WRITE_2_SUB=>
		ESTADO <= WRITE_2_EN_SUB;
		
		WHEN WRITE_2_EN_SUB =>
		ESTADO<= SUB_MENU_Y;

		
		WHEN WRITE_RXR3_SUB=>
		ESTADO<=WRITE_RXR3_ADDRESS1_SUB;
		
		WHEN WRITE_RXR3_ADDRESS1_SUB=>
		ESTADO<= WRITE_RXR3_1_SUB;
		
		WHEN WRITE_RXR3_1_SUB=>
		ESTADO<= WRITE_RXR3_1_EN_SUB;
		
		WHEN WRITE_RXR3_1_EN_SUB=>
		ESTADO<= WRITE_RXR3_ADDRESS2_SUB;
		
		WHEN WRITE_RXR3_ADDRESS2_SUB=>
		ESTADO<= WRITE_RXR3_ADDRESS2_EN_SUB;
		
		WHEN WRITE_RXR3_ADDRESS2_EN_SUB=>
		ESTADO<= WRITE_3_SUB;
		
		WHEN WRITE_3_SUB=>
		ESTADO <= WRITE_3_EN_SUB;
		
		WHEN WRITE_3_EN_SUB =>
		ESTADO<= SUB_MENU_Y;
		
		WHEN WRITE_RX_SUB=>
		ESTADO<=WRITE_RX_ADDRESS1_SUB;
		
		WHEN WRITE_RX_ADDRESS1_SUB=>
		ESTADO<= WRITE_RX_1_SUB;
		
		WHEN WRITE_RX_1_SUB=>
		ESTADO<= WRITE_RX_1_EN_SUB;
		
		WHEN WRITE_RX_1_EN_SUB=>
		ESTADO<= WRITE_RX_ADDRESS2_SUB;
		
		WHEN WRITE_RX_ADDRESS2_SUB=>
		ESTADO<= WRITE_RX_ADDRESS2_EN_SUB;
		
		WHEN WRITE_RX_ADDRESS2_EN_SUB=>
		ESTADO<= WRITE_x_SUB;
		
		WHEN WRITE_x_SUB=>
		ESTADO <= WRITE_x_EN_SUB;
		
		WHEN WRITE_x_EN_SUB =>
		ESTADO<= SUB_MENU_Y;
		
		
		
		

		WHEN WRITE_RYR1_SUB=>
		ESTADO<=WRITE_RYR1_ADDRESS1_SUB;
		
		WHEN WRITE_RYR1_ADDRESS1_SUB=>
		ESTADO<= WRITE_1Y_SUB;
		
		WHEN WRITE_1Y_SUB=>
		ESTADO <= WRITE_1Y_EN_SUB;
		
		WHEN WRITE_1Y_EN_SUB =>
		ESTADO<= SUB_MENU_X;

		
		WHEN WRITE_RYR2_SUB=>
		ESTADO<=WRITE_RYR2_ADDRESS1_SUB;
		
		WHEN WRITE_RYR2_ADDRESS1_SUB=>
		ESTADO<= WRITE_2Y_SUB;
		
		WHEN WRITE_2Y_SUB=>
		ESTADO <= WRITE_2Y_EN_SUB;
		
		WHEN WRITE_2Y_EN_SUB =>
		ESTADO<= SUB_MENU_X;

		
		
		WHEN WRITE_RYR3_SUB=>
		ESTADO<=WRITE_RYR3_ADDRESS1_SUB;
		
		WHEN WRITE_RYR3_ADDRESS1_SUB=>
		ESTADO<= WRITE_3Y_SUB;
		
		WHEN WRITE_3Y_SUB=>
		ESTADO <= WRITE_3Y_EN_SUB;
		
		WHEN WRITE_3Y_EN_SUB =>
		ESTADO<= SUB_MENU_X;
		
		
		
		WHEN WRITE_RY_SUB=>
		ESTADO<=WRITE_RY_ADDRESS1_SUB;
		
		WHEN WRITE_RY_ADDRESS1_SUB=>
		ESTADO<= WRITE_Y_SUB;
		
		WHEN WRITE_Y_SUB=>
		ESTADO <= WRITE_Y_EN_SUB;
		
		WHEN WRITE_Y_EN_SUB =>
		ESTADO<= SUB_MENU_X;

-------------------------------------------------------------------------
---------------------------------------------------------------
		
		
		WHEN WRITE_RXR1_AND=>
		ESTADO<=WRITE_RXR1_ADDRESS1_AND;
		
		WHEN WRITE_RXR1_ADDRESS1_AND=>
		ESTADO<= WRITE_RXR1_1_AND;
		
		WHEN WRITE_RXR1_1_AND=>
		ESTADO<= WRITE_RXR1_1_EN_AND;
		
		WHEN WRITE_RXR1_1_EN_AND=>
		ESTADO<= WRITE_RXR1_ADDRESS2_AND;
		
		WHEN WRITE_RXR1_ADDRESS2_AND=>
		ESTADO<= WRITE_RXR1_ADDRESS2_EN_AND;
		
		WHEN WRITE_RXR1_ADDRESS2_EN_AND=>
		ESTADO<= WRITE_1_AND;
		
		WHEN WRITE_1_AND=>
		ESTADO <= WRITE_1_EN_AND;
		
		WHEN WRITE_1_EN_AND =>
		ESTADO<= AND_MENU_Y;
		
		
		WHEN WRITE_RXR2_AND=>
		ESTADO<=WRITE_RXR2_ADDRESS1_AND;
		
		WHEN WRITE_RXR2_ADDRESS1_AND=>
		ESTADO<= WRITE_RXR2_1_AND;
		
		WHEN WRITE_RXR2_1_AND=>
		ESTADO<= WRITE_RXR2_1_EN_AND;
		
		WHEN WRITE_RXR2_1_EN_AND=>
		ESTADO<= WRITE_RXR2_ADDRESS2_AND;
		
		WHEN WRITE_RXR2_ADDRESS2_AND=>
		ESTADO<= WRITE_RXR2_ADDRESS2_EN_AND;
		
		WHEN WRITE_RXR2_ADDRESS2_EN_AND=>
		ESTADO<= WRITE_2_AND;
		
		WHEN WRITE_2_AND=>
		ESTADO <= WRITE_2_EN_AND;
		
		WHEN WRITE_2_EN_AND =>
		ESTADO<= AND_MENU_Y;

		
		WHEN WRITE_RXR3_AND=>
		ESTADO<=WRITE_RXR3_ADDRESS1_AND;
		
		WHEN WRITE_RXR3_ADDRESS1_AND=>
		ESTADO<= WRITE_RXR3_1_AND;
		
		WHEN WRITE_RXR3_1_AND=>
		ESTADO<= WRITE_RXR3_1_EN_AND;
		
		WHEN WRITE_RXR3_1_EN_AND=>
		ESTADO<= WRITE_RXR3_ADDRESS2_AND;
		
		WHEN WRITE_RXR3_ADDRESS2_AND=>
		ESTADO<= WRITE_RXR3_ADDRESS2_EN_AND;
		
		WHEN WRITE_RXR3_ADDRESS2_EN_AND=>
		ESTADO<= WRITE_3_AND;
		
		WHEN WRITE_3_AND=>
		ESTADO <= WRITE_3_EN_AND;
		
		WHEN WRITE_3_EN_AND =>
		ESTADO<= AND_MENU_Y;
		
		WHEN WRITE_RX_AND=>
		ESTADO<=WRITE_RX_ADDRESS1_AND;
		
		WHEN WRITE_RX_ADDRESS1_AND=>
		ESTADO<= WRITE_RX_1_AND;
		
		WHEN WRITE_RX_1_AND=>
		ESTADO<= WRITE_RX_1_EN_AND;
		
		WHEN WRITE_RX_1_EN_AND=>
		ESTADO<= WRITE_RX_ADDRESS2_AND;
		
		WHEN WRITE_RX_ADDRESS2_AND=>
		ESTADO<= WRITE_RX_ADDRESS2_EN_AND;
		
		WHEN WRITE_RX_ADDRESS2_EN_AND=>
		ESTADO<= WRITE_x_AND;
		
		WHEN WRITE_x_AND=>
		ESTADO <= WRITE_x_EN_AND;
		
		WHEN WRITE_x_EN_AND =>
		ESTADO<= AND_MENU_Y;
		
		
		
		

		WHEN WRITE_RYR1_AND=>
		ESTADO<=WRITE_RYR1_ADDRESS1_AND;
		
		WHEN WRITE_RYR1_ADDRESS1_AND=>
		ESTADO<= WRITE_1Y_AND;
		
		WHEN WRITE_1Y_AND=>
		ESTADO <= WRITE_1Y_EN_AND;
		
		WHEN WRITE_1Y_EN_AND =>
		ESTADO<= AND_MENU_X;

		
		WHEN WRITE_RYR2_AND=>
		ESTADO<=WRITE_RYR2_ADDRESS1_AND;
		
		WHEN WRITE_RYR2_ADDRESS1_AND=>
		ESTADO<= WRITE_2Y_AND;
		
		WHEN WRITE_2Y_AND=>
		ESTADO <= WRITE_2Y_EN_AND;
		
		WHEN WRITE_2Y_EN_AND =>
		ESTADO<= AND_MENU_X;

		
		
		WHEN WRITE_RYR3_AND=>
		ESTADO<=WRITE_RYR3_ADDRESS1_AND;
		
		WHEN WRITE_RYR3_ADDRESS1_AND=>
		ESTADO<= WRITE_3Y_AND;
		
		WHEN WRITE_3Y_AND=>
		ESTADO <= WRITE_3Y_EN_AND;
		
		WHEN WRITE_3Y_EN_AND =>
		ESTADO<= AND_MENU_X;
		
		
		
		WHEN WRITE_RY_AND=>
		ESTADO<=WRITE_RY_ADDRESS1_AND;
		
		WHEN WRITE_RY_ADDRESS1_AND=>
		ESTADO<= WRITE_Y_AND;
		
		WHEN WRITE_Y_AND=>
		ESTADO <= WRITE_Y_EN_AND;
		
		WHEN WRITE_Y_EN_AND =>
		ESTADO<= AND_MENU_X;

-------------------------------------------------------------------------
---------------------------------------------------------------
		
		
		WHEN WRITE_RXR1_NOT=>
		ESTADO<=WRITE_RXR1_ADDRESS1_NOT;
		
		WHEN WRITE_RXR1_ADDRESS1_NOT=>
		ESTADO<= WRITE_RXR1_1_NOT;
		
		WHEN WRITE_RXR1_1_NOT=>
		ESTADO<= WRITE_RXR1_1_EN_NOT;
		
		WHEN WRITE_RXR1_1_EN_NOT=>
		ESTADO<= NOT_MENU_Y;
		
		
		WHEN WRITE_RXR2_NOT=>
		ESTADO<=WRITE_RXR2_ADDRESS1_NOT;
		
		WHEN WRITE_RXR2_ADDRESS1_NOT=>
		ESTADO<= WRITE_RXR2_1_NOT;
		
		WHEN WRITE_RXR2_1_NOT=>
		ESTADO<= WRITE_RXR2_1_EN_NOT;
		
		WHEN WRITE_RXR2_1_EN_NOT=>
		ESTADO<= NOT_MENU_Y;
		

		
		WHEN WRITE_RXR3_NOT=>
		ESTADO<=WRITE_RXR3_ADDRESS1_NOT;
		
		WHEN WRITE_RXR3_ADDRESS1_NOT=>
		ESTADO<= WRITE_RXR3_1_NOT;
		
		WHEN WRITE_RXR3_1_NOT=>
		ESTADO<= WRITE_RXR3_1_EN_NOT;
		
		WHEN WRITE_RXR3_1_EN_NOT=>
		ESTADO<= NOT_MENU_Y;
		
		
		WHEN WRITE_RX_NOT=>
		ESTADO<=WRITE_RX_ADDRESS1_NOT;
		
		WHEN WRITE_RX_ADDRESS1_NOT=>
		ESTADO<= WRITE_RX_1_NOT;
		
		WHEN WRITE_RX_1_NOT=>
		ESTADO<= WRITE_RX_1_EN_NOT;
		
		WHEN WRITE_RX_1_EN_NOT=>
		ESTADO<= NOT_MENU_Y;
		
		
		

		WHEN WRITE_RYR1_NOT=>
		ESTADO<=WRITE_RYR1_ADDRESS1_NOT;
		
		WHEN WRITE_RYR1_ADDRESS1_NOT=>
		ESTADO<= WRITE_RYR1_1_NOT;
		
		WHEN WRITE_RYR1_1_NOT=>
		ESTADO <= WRITE_RYR1_1_EN_NOT;
		
		WHEN WRITE_RYR1_1_EN_NOT =>
		ESTADO<= NOT_MENU_X;

		
		WHEN WRITE_RYR2_NOT=>
		ESTADO<=WRITE_RYR2_ADDRESS1_NOT;
		
		WHEN WRITE_RYR2_ADDRESS1_NOT=>
		ESTADO<= WRITE_RYR2_1_NOT;
		
		WHEN WRITE_RYR2_1_NOT=>
		ESTADO <= WRITE_RYR2_1_EN_NOT;
		
		WHEN WRITE_RYR2_1_EN_NOT =>
		ESTADO<= NOT_MENU_X;

		
		
		WHEN WRITE_RYR3_NOT=>
		ESTADO<=WRITE_RYR3_ADDRESS1_NOT;
		
		WHEN WRITE_RYR3_ADDRESS1_NOT=>
		ESTADO<= WRITE_RYR3_1_NOT;
		
		WHEN WRITE_RYR3_1_NOT=>
		ESTADO <= WRITE_RYR3_1_EN_NOT;
		
		WHEN WRITE_RYR3_1_EN_NOT=>
		ESTADO<= NOT_MENU_X;
		
		
		
		WHEN WRITE_RY_NOT=>
		ESTADO<=WRITE_RY_ADDRESS1_NOT;
		
		WHEN WRITE_RY_ADDRESS1_NOT=>
		ESTADO<= WRITE_RY_1_NOT;
		
		WHEN WRITE_RY_1_NOT=>
		ESTADO <= WRITE_RY_1_EN_NOT;
		
		WHEN WRITE_RY_1_EN_NOT =>
		ESTADO<= NOT_MENU_X;

-------------------------------------------------------------------------
-------------------------------------------------------------------------		
		
		WHEN WRITE_RXR1_SWAP=>
		ESTADO<=WRITE_RXR1_ADDRESS1_SWAP;
		
		WHEN WRITE_RXR1_ADDRESS1_SWAP=>
		ESTADO<= WRITE_RXR1_1_SWAP;
		
		WHEN WRITE_RXR1_1_SWAP=>
		ESTADO<= WRITE_RXR1_1_EN_SWAP;
		
		WHEN WRITE_RXR1_1_EN_SWAP=>
		ESTADO<= SWAP_MENU_Y;
		
		
		WHEN WRITE_RXR2_SWAP=>
		ESTADO<=WRITE_RXR2_ADDRESS1_SWAP;
		
		WHEN WRITE_RXR2_ADDRESS1_SWAP=>
		ESTADO<= WRITE_RXR2_1_SWAP;
		
		WHEN WRITE_RXR2_1_SWAP=>
		ESTADO<= WRITE_RXR2_1_EN_SWAP;
		
		WHEN WRITE_RXR2_1_EN_SWAP=>
		ESTADO<= SWAP_MENU_Y;
		

		
		WHEN WRITE_RXR3_SWAP=>
		ESTADO<=WRITE_RXR3_ADDRESS1_SWAP;
		
		WHEN WRITE_RXR3_ADDRESS1_SWAP=>
		ESTADO<= WRITE_RXR3_1_SWAP;
		
		WHEN WRITE_RXR3_1_SWAP=>
		ESTADO<= WRITE_RXR3_1_EN_SWAP;
		
		WHEN WRITE_RXR3_1_EN_SWAP=>
		ESTADO<= SWAP_MENU_Y;
		
		
		WHEN WRITE_RX_SWAP=>
		ESTADO<=WRITE_RX_ADDRESS1_SWAP;
		
		WHEN WRITE_RX_ADDRESS1_SWAP=>
		ESTADO<= WRITE_RX_1_SWAP;
		
		WHEN WRITE_RX_1_SWAP=>
		ESTADO<= WRITE_RX_1_EN_SWAP;
		
		WHEN WRITE_RX_1_EN_SWAP=>
		ESTADO<= SWAP_MENU_Y;
		
		
		

		WHEN WRITE_RYR1_SWAP=>
		ESTADO<=WRITE_RYR1_ADDRESS1_SWAP;
		
		WHEN WRITE_RYR1_ADDRESS1_SWAP=>
		ESTADO<= WRITE_RYR1_1_SWAP;
		
		WHEN WRITE_RYR1_1_SWAP=>
		ESTADO <= WRITE_RYR1_1_EN_SWAP;
		
		WHEN WRITE_RYR1_1_EN_SWAP =>
		ESTADO<= SWAP_MENU_X;

		
		WHEN WRITE_RYR2_SWAP=>
		ESTADO<=WRITE_RYR2_ADDRESS1_SWAP;
		
		WHEN WRITE_RYR2_ADDRESS1_SWAP=>
		ESTADO<= WRITE_RYR2_1_SWAP;
		
		WHEN WRITE_RYR2_1_SWAP=>
		ESTADO <= WRITE_RYR2_1_EN_SWAP;
		
		WHEN WRITE_RYR2_1_EN_SWAP=>
		ESTADO<= SWAP_MENU_X;

		
		
		WHEN WRITE_RYR3_SWAP=>
		ESTADO<=WRITE_RYR3_ADDRESS1_SWAP;
		
		WHEN WRITE_RYR3_ADDRESS1_SWAP=>
		ESTADO<= WRITE_RYR3_1_SWAP;
		
		WHEN WRITE_RYR3_1_SWAP=>
		ESTADO <= WRITE_RYR3_1_EN_SWAP;
		
		WHEN WRITE_RYR3_1_EN_SWAP=>
		ESTADO<= SWAP_MENU_X;
		
		
		
		WHEN WRITE_RY_SWAP=>
		ESTADO<=WRITE_RY_ADDRESS1_SWAP;
		
		WHEN WRITE_RY_ADDRESS1_SWAP=>
		ESTADO<= WRITE_RY_1_SWAP;
		
		WHEN WRITE_RY_1_SWAP=>
		ESTADO <= WRITE_RY_1_EN_SWAP;
		
		WHEN WRITE_RY_1_EN_SWAP=>
		ESTADO<= SWAP_MENU_X;


---------------------------------------------------------------
---------------------------------------------------------------
		
		WHEN WRITE_RXR1_OR=>
		ESTADO<=WRITE_RXR1_ADDRESS1_OR;
		
		WHEN WRITE_RXR1_ADDRESS1_OR=>
		ESTADO<= WRITE_RXR1_1_OR;
		
		WHEN WRITE_RXR1_1_OR=>
		ESTADO<= WRITE_RXR1_1_EN_OR;
		
		WHEN WRITE_RXR1_1_EN_OR=>
		ESTADO<= WRITE_RXR1_ADDRESS2_OR;
		
		WHEN WRITE_RXR1_ADDRESS2_OR=>
		ESTADO<= WRITE_RXR1_ADDRESS2_EN_OR;
		
		WHEN WRITE_RXR1_ADDRESS2_EN_OR=>
		ESTADO<= WRITE_1_OR;
		
		WHEN WRITE_1_OR=>
		ESTADO <= WRITE_1_EN_OR;
		
		WHEN WRITE_1_EN_OR =>
		ESTADO<= OR_MENU_Y;
		
		
		WHEN WRITE_RXR2_OR=>
		ESTADO<=WRITE_RXR2_ADDRESS1_OR;
		
		WHEN WRITE_RXR2_ADDRESS1_OR=>
		ESTADO<= WRITE_RXR2_1_OR;
		
		WHEN WRITE_RXR2_1_OR=>
		ESTADO<= WRITE_RXR2_1_EN_OR;
		
		WHEN WRITE_RXR2_1_EN_OR=>
		ESTADO<= WRITE_RXR2_ADDRESS2_OR;
		
		WHEN WRITE_RXR2_ADDRESS2_OR=>
		ESTADO<= WRITE_RXR2_ADDRESS2_EN_OR;
		
		WHEN WRITE_RXR2_ADDRESS2_EN_OR=>
		ESTADO<= WRITE_2_OR;
		
		WHEN WRITE_2_OR=>
		ESTADO <= WRITE_2_EN_OR;
		
		WHEN WRITE_2_EN_OR =>
		ESTADO<= OR_MENU_Y;

		
		WHEN WRITE_RXR3_OR=>
		ESTADO<=WRITE_RXR3_ADDRESS1_OR;
		
		WHEN WRITE_RXR3_ADDRESS1_OR=>
		ESTADO<= WRITE_RXR3_1_OR;
		
		WHEN WRITE_RXR3_1_OR=>
		ESTADO<= WRITE_RXR3_1_EN_OR;
		
		WHEN WRITE_RXR3_1_EN_OR=>
		ESTADO<= WRITE_RXR3_ADDRESS2_OR;
		
		WHEN WRITE_RXR3_ADDRESS2_OR=>
		ESTADO<= WRITE_RXR3_ADDRESS2_EN_OR;
		
		WHEN WRITE_RXR3_ADDRESS2_EN_OR=>
		ESTADO<= WRITE_3_OR;
		
		WHEN WRITE_3_OR=>
		ESTADO <= WRITE_3_EN_OR;
		
		WHEN WRITE_3_EN_OR =>
		ESTADO<= OR_MENU_Y;
		
		WHEN WRITE_RX_OR=>
		ESTADO<=WRITE_RX_ADDRESS1_OR;
		
		WHEN WRITE_RX_ADDRESS1_OR=>
		ESTADO<= WRITE_RX_1_OR;
		
		WHEN WRITE_RX_1_OR=>
		ESTADO<= WRITE_RX_1_EN_OR;
		
		WHEN WRITE_RX_1_EN_OR=>
		ESTADO<= WRITE_RX_ADDRESS2_OR;
		
		WHEN WRITE_RX_ADDRESS2_OR=>
		ESTADO<= WRITE_RX_ADDRESS2_EN_OR;
		
		WHEN WRITE_RX_ADDRESS2_EN_OR=>
		ESTADO<= WRITE_x_OR;
		
		WHEN WRITE_x_OR=>
		ESTADO <= WRITE_x_EN_OR;
		
		WHEN WRITE_x_EN_OR =>
		ESTADO<= OR_MENU_Y;
		
		
		
		

		WHEN WRITE_RYR1_OR=>
		ESTADO<=WRITE_RYR1_ADDRESS1_OR;
		
		WHEN WRITE_RYR1_ADDRESS1_OR=>
		ESTADO<= WRITE_1Y_OR;
		
		WHEN WRITE_1Y_OR=>
		ESTADO <= WRITE_1Y_EN_OR;
		
		WHEN WRITE_1Y_EN_OR =>
		ESTADO<= OR_MENU_X;

		
		WHEN WRITE_RYR2_OR=>
		ESTADO<=WRITE_RYR2_ADDRESS1_OR;
		
		WHEN WRITE_RYR2_ADDRESS1_OR=>
		ESTADO<= WRITE_2Y_OR;
		
		WHEN WRITE_2Y_OR=>
		ESTADO <= WRITE_2Y_EN_OR;
		
		WHEN WRITE_2Y_EN_OR =>
		ESTADO<= OR_MENU_X;

		
		
		WHEN WRITE_RYR3_OR=>
		ESTADO<=WRITE_RYR3_ADDRESS1_OR;
		
		WHEN WRITE_RYR3_ADDRESS1_OR=>
		ESTADO<= WRITE_3Y_OR;
		
		WHEN WRITE_3Y_OR=>
		ESTADO <= WRITE_3Y_EN_OR;
		
		WHEN WRITE_3Y_EN_OR =>
		ESTADO<= OR_MENU_X;
		
		
		
		WHEN WRITE_RY_OR=>
		ESTADO<=WRITE_RY_ADDRESS1_OR;
		
		WHEN WRITE_RY_ADDRESS1_OR=>
		ESTADO<= WRITE_Y_OR;
		
		WHEN WRITE_Y_OR=>
		ESTADO <= WRITE_Y_EN_OR;
		
		WHEN WRITE_Y_EN_OR =>
		ESTADO<= OR_MENU_X;

-------------------------------------------------------------------------
---------------------------------------------------------------
		
		
		WHEN WRITE_RXR1_MUL=>
		ESTADO<=WRITE_RXR1_ADDRESS1_MUL;
		
		WHEN WRITE_RXR1_ADDRESS1_MUL=>
		ESTADO<= WRITE_RXR1_1_MUL;
		
		WHEN WRITE_RXR1_1_MUL=>
		ESTADO<= WRITE_RXR1_1_EN_MUL;
		
		WHEN WRITE_RXR1_1_EN_MUL=>
		ESTADO<= WRITE_RXR1_ADDRESS2_MUL;
		
		WHEN WRITE_RXR1_ADDRESS2_MUL=>
		ESTADO<= WRITE_RXR1_ADDRESS2_EN_MUL;
		
		WHEN WRITE_RXR1_ADDRESS2_EN_MUL=>
		ESTADO<= WRITE_1_MUL;
		
		WHEN WRITE_1_MUL=>
		ESTADO <= WRITE_1_EN_MUL;
		
		WHEN WRITE_1_EN_MUL =>
		ESTADO<= MUL_MENU_Y;

		
		WHEN WRITE_RXR2_MUL=>
		ESTADO<=WRITE_RXR2_ADDRESS1_MUL;
		
		WHEN WRITE_RXR2_ADDRESS1_MUL=>
		ESTADO<= WRITE_RXR2_1_MUL;
		
		WHEN WRITE_RXR2_1_MUL=>
		ESTADO<= WRITE_RXR2_1_EN_MUL;
		
		WHEN WRITE_RXR2_1_EN_MUL=>
		ESTADO<= WRITE_RXR2_ADDRESS2_MUL;
		
		WHEN WRITE_RXR2_ADDRESS2_MUL=>
		ESTADO<= WRITE_RXR2_ADDRESS2_EN_MUL;
		
		WHEN WRITE_RXR2_ADDRESS2_EN_MUL=>
		ESTADO<= WRITE_2_MUL;
		
		WHEN WRITE_2_MUL=>
		ESTADO <= WRITE_2_EN_MUL;
		
		WHEN WRITE_2_EN_MUL =>
		ESTADO<= MUL_MENU_Y;

		
		WHEN WRITE_RXR3_MUL=>
		ESTADO<=WRITE_RXR3_ADDRESS1_MUL;
		
		WHEN WRITE_RXR3_ADDRESS1_MUL=>
		ESTADO<= WRITE_RXR3_1_MUL;
		
		WHEN WRITE_RXR3_1_MUL=>
		ESTADO<= WRITE_RXR3_1_EN_MUL;
		
		WHEN WRITE_RXR3_1_EN_MUL=>
		ESTADO<= WRITE_RXR3_ADDRESS2_MUL;
		
		WHEN WRITE_RXR3_ADDRESS2_MUL=>
		ESTADO<= WRITE_RXR3_ADDRESS2_EN_MUL;
		
		WHEN WRITE_RXR3_ADDRESS2_EN_MUL=>
		ESTADO<= WRITE_3_MUL;
		
		WHEN WRITE_3_MUL=>
		ESTADO <= WRITE_3_EN_MUL;
		
		WHEN WRITE_3_EN_MUL =>
		ESTADO<= MUL_MENU_Y;
		
		
		WHEN WRITE_RX_MUL=>
		ESTADO<=WRITE_RX_ADDRESS1_MUL;
		
		WHEN WRITE_RX_ADDRESS1_MUL=>
		ESTADO<= WRITE_RX_1_MUL;
		
		WHEN WRITE_RX_1_MUL=>
		ESTADO<= WRITE_RX_1_EN_MUL;
		
		WHEN WRITE_RX_1_EN_MUL=>
		ESTADO<= WRITE_RX_ADDRESS2_MUL;
		
		WHEN WRITE_RX_ADDRESS2_MUL=>
		ESTADO<= WRITE_RX_ADDRESS2_EN_MUL;
		
		WHEN WRITE_RX_ADDRESS2_EN_MUL=>
		ESTADO<= WRITE_x_MUL;
		
		WHEN WRITE_x_MUL=>
		ESTADO <= WRITE_x_EN_MUL;
		
		WHEN WRITE_x_EN_MUL =>
		ESTADO<= MUL_MENU_Y;
		
		
		
		

		WHEN WRITE_RYR1_MUL=>
		ESTADO<=WRITE_RYR1_ADDRESS1_MUL;
		
		WHEN WRITE_RYR1_ADDRESS1_MUL=>
		ESTADO<= WRITE_1Y_MUL;
		
		WHEN WRITE_1Y_MUL=>
		ESTADO <= WRITE_1Y_EN_MUL;
		
		WHEN WRITE_1Y_EN_MUL =>
		ESTADO<= MUL_MENU_X;

		
		WHEN WRITE_RYR2_MUL=>
		ESTADO<=WRITE_RYR2_ADDRESS1_MUL;
		
		WHEN WRITE_RYR2_ADDRESS1_MUL=>
		ESTADO<= WRITE_2Y_MUL;
		
		WHEN WRITE_2Y_MUL=>
		ESTADO <= WRITE_2Y_EN_MUL;
		
		WHEN WRITE_2Y_EN_MUL =>
		ESTADO<= MUL_MENU_X;

		
		
		WHEN WRITE_RYR3_MUL=>
		ESTADO<=WRITE_RYR3_ADDRESS1_MUL;
		
		WHEN WRITE_RYR3_ADDRESS1_MUL=>
		ESTADO<= WRITE_3Y_MUL;
		
		WHEN WRITE_3Y_MUL=>
		ESTADO <= WRITE_3Y_EN_MUL;
		
		WHEN WRITE_3Y_EN_MUL =>
		ESTADO<= MUL_MENU_X;
		
		
		
		WHEN WRITE_RY_MUL=>
		ESTADO<=WRITE_RY_ADDRESS1_MUL;
		
		WHEN WRITE_RY_ADDRESS1_MUL=>
		ESTADO<= WRITE_Y_MUL;
		
		WHEN WRITE_Y_MUL=>
		ESTADO <= WRITE_Y_EN_MUL;
		
		WHEN WRITE_Y_EN_MUL =>
		ESTADO<= MUL_MENU_X;

-------------------------------------------------------------------------
-------------------------------------------------------------------------
		WHEN WRITE_RYR1_LOAD=>
		ESTADO<=WRITE_RYR1_ADDRESS1_LOAD;
		
		WHEN WRITE_RYR1_ADDRESS1_LOAD=>
		ESTADO<= WRITE_1Y_LOAD;
		
		WHEN WRITE_1Y_LOAD=>
		ESTADO <= WRITE_1Y_EN_LOAD;
		
		WHEN WRITE_1Y_EN_LOAD =>
		ESTADO<= LOAD_MENU_Y;

		
		WHEN WRITE_RYR2_LOAD=>
		ESTADO<=WRITE_RYR2_ADDRESS1_LOAD;
		
		WHEN WRITE_RYR2_ADDRESS1_LOAD=>
		ESTADO<= WRITE_2Y_LOAD;
		
		WHEN WRITE_2Y_LOAD=>
		ESTADO <= WRITE_2Y_EN_LOAD;
		
		WHEN WRITE_2Y_EN_LOAD =>
		ESTADO<= LOAD_MENU_Y;

		
		
		WHEN WRITE_RYR3_LOAD=>
		ESTADO<=WRITE_RYR3_ADDRESS1_LOAD;
		
		WHEN WRITE_RYR3_ADDRESS1_LOAD=>
		ESTADO<= WRITE_3Y_LOAD;
		
		WHEN WRITE_3Y_LOAD=>
		ESTADO <= WRITE_3Y_EN_LOAD;
		
		WHEN WRITE_3Y_EN_LOAD =>
		ESTADO<= LOAD_MENU_Y;
		
		
		
		WHEN WRITE_RY_LOAD=>
		ESTADO<=WRITE_RY_ADDRESS1_LOAD;
		
		WHEN WRITE_RY_ADDRESS1_LOAD=>
		ESTADO<= WRITE_Y_LOAD;
		
		WHEN WRITE_Y_LOAD=>
		ESTADO <= WRITE_Y_EN_LOAD;
		
		WHEN WRITE_Y_EN_LOAD =>
		ESTADO<= LOAD_MENU_Y;
------------------------------------------------------------------------
------------------------------------------------------------------------
		
		WHEN WRITE_RXR1_COMP=>
		ESTADO<=WRITE_RXR1_ADDRESS1_COMP;
		
		WHEN WRITE_RXR1_ADDRESS1_COMP=>
		ESTADO<= WRITE_RXR1_1_COMP;
		
		WHEN WRITE_RXR1_1_COMP=>
		ESTADO<= WRITE_RXR1_1_EN_COMP;
		
		WHEN WRITE_RXR1_1_EN_COMP=>
		ESTADO<= COMP_MENU_Y;
		
		
		WHEN WRITE_RXR2_COMP=>
		ESTADO<=WRITE_RXR2_ADDRESS1_COMP;
		
		WHEN WRITE_RXR2_ADDRESS1_COMP=>
		ESTADO<= WRITE_RXR2_1_COMP;
		
		WHEN WRITE_RXR2_1_COMP=>
		ESTADO<= WRITE_RXR2_1_EN_COMP;
		
		WHEN WRITE_RXR2_1_EN_COMP=>
		ESTADO<= COMP_MENU_Y;
		

		
		WHEN WRITE_RXR3_COMP=>
		ESTADO<=WRITE_RXR3_ADDRESS1_COMP;
		
		WHEN WRITE_RXR3_ADDRESS1_COMP=>
		ESTADO<= WRITE_RXR3_1_COMP;
		
		WHEN WRITE_RXR3_1_COMP=>
		ESTADO<= WRITE_RXR3_1_EN_COMP;
		
		WHEN WRITE_RXR3_1_EN_COMP=>
		ESTADO<= COMP_MENU_Y;
		
		
		WHEN WRITE_RX_COMP=>
		ESTADO<=WRITE_RX_ADDRESS1_COMP;
		
		WHEN WRITE_RX_ADDRESS1_COMP=>
		ESTADO<= WRITE_RX_1_COMP;
		
		WHEN WRITE_RX_1_COMP=>
		ESTADO<= WRITE_RX_1_EN_COMP;
		
		WHEN WRITE_RX_1_EN_COMP=>
		ESTADO<= COMP_MENU_Y;
		
		
		

		WHEN WRITE_RYR1_COMP=>
		ESTADO<=WRITE_RYR1_ADDRESS1_COMP;
		
		WHEN WRITE_RYR1_ADDRESS1_COMP=>
		ESTADO<= WRITE_RYR1_1_COMP;
		
		WHEN WRITE_RYR1_1_COMP=>
		ESTADO <= WRITE_RYR1_1_EN_COMP;
		
		WHEN WRITE_RYR1_1_EN_COMP=>
		ESTADO<= COMP_MENU_OPERATOR;

		
		WHEN WRITE_RYR2_COMP=>
		ESTADO<=WRITE_RYR2_ADDRESS1_COMP;
		
		WHEN WRITE_RYR2_ADDRESS1_COMP=>
		ESTADO<= WRITE_RYR2_1_COMP;
		
		WHEN WRITE_RYR2_1_COMP=>
		ESTADO <= WRITE_RYR2_1_EN_COMP;
		
		WHEN WRITE_RYR2_1_EN_COMP=>
		ESTADO<= COMP_MENU_OPERATOR;

		
		
		WHEN WRITE_RYR3_COMP=>
		ESTADO<=WRITE_RYR3_ADDRESS1_COMP;
		
		WHEN WRITE_RYR3_ADDRESS1_COMP=>
		ESTADO<= WRITE_RYR3_1_COMP;
		
		WHEN WRITE_RYR3_1_COMP=>
		ESTADO <= WRITE_RYR3_1_EN_COMP;
		
		WHEN WRITE_RYR3_1_EN_COMP=>
		ESTADO<= COMP_MENU_OPERATOR;
		
		
		
		WHEN WRITE_RY_COMP=>
		ESTADO<=WRITE_RY_ADDRESS1_COMP;
		
		WHEN WRITE_RY_ADDRESS1_COMP=>
		ESTADO<= WRITE_RY_1_COMP;
		
		WHEN WRITE_RY_1_COMP=>
		ESTADO <= WRITE_RY_1_EN_COMP;
		
		WHEN WRITE_RY_1_EN_COMP=>
		ESTADO<= COMP_MENU_OPERATOR;
		
		
		-- Note que no caso da comparação temos algumas etapas a mais de interpretação referentes aos sinais
		-- de EQU,GRT e LST, que também são mostrados no display LCD
		
		WHEN COMP_ADDRESS_OPERATOR=>
		ESTADO<= COMP_ADDRESS_OPERATOR_EN;
		
		WHEN COMP_ADDRESS_OPERATOR_EN=>
		IF ENABLE = '0' THEN
		ESTADO<= COMP_WAIT;
		ELSIF (ENABLE = '1') AND (GRT = '1') THEN
		ESTADO<= COMP_MAIOR;
	
		ELSIF (ENABLE = '1') AND (LST = '1') THEN
		ESTADO<= COMP_MENOR;
		
		ELSIF (ENABLE = '1') AND (EQU = '1') THEN
		ESTADO<= COMP_IGUAL;
		END IF;
		
		
		WHEN COMP_WAIT =>
		ESTADO <= COMP_WAIT_EN;
		
		WHEN COMP_WAIT_EN =>
		ESTADO <= COMP_MENU_X;
		
		
		WHEN COMP_MAIOR =>
		ESTADO <= COMP_MAIOR_EN;
		
		WHEN COMP_MAIOR_EN =>
		ESTADO <= COMP_MENU_X;
		
		
		WHEN COMP_MENOR =>
		ESTADO <= COMP_MENOR_EN;
		
		WHEN COMP_MENOR_EN =>
		ESTADO <= COMP_MENU_X;
		
		
		WHEN COMP_IGUAL =>
		ESTADO <= COMP_IGUAL_EN;
		
		WHEN COMP_IGUAL_EN =>
		ESTADO <= COMP_MENU_X;
-------------------------------------------------------------------------

		WHEN OTHERS=>
		NULL;
		END CASE;
	END IF;
END PROCESS;

-- O case abaixo é responsável por realizar a manipulação dos sinais referentes em cada estado
PROCESS (ESTADO)
BEGIN
	CASE ESTADO IS
		WHEN IDLE_CLEAR1 =>
				LCD_DATA <= CDG_iniciacao(conteiro);
				LCD_EN <= '1';
				LCD_RW <= '0';
				LCD_RS <= '0';
				
		WHEN IDLE_CLEAR2 =>
				LCD_EN <= '0';
				LCD_RW <= '0';
				LCD_RS <= '0';
			
		WHEN IDLE =>
				LCD_EN <= '0';
				LCD_RW <= '0';
				LCD_RS <= '0';
			
		WHEN LINHA1_ADDRESS_SET=>
				LCD_DATA <="10000000";
				LCD_EN <= '1';
				LCD_RW <= '0';
				LCD_RS <= '0';
				
		WHEN LINHA1_ADDRESS_EN=>
				LCD_EN <= '0';
				LCD_RW <= '0';
				LCD_RS <= '0';

		WHEN LINHA2_ADDRESS_SET=>
				LCD_DATA <="11000000";
				LCD_EN <= '1';
				LCD_RW <= '0';
				LCD_RS <= '0';
				
		WHEN LINHA2_ADDRESS_EN=>
				LCD_EN <= '0';
				LCD_RW <= '0';
				LCD_RS <= '0';
				
		WHEN LOAD_MSG =>
				LCD_DATA <= Linha_LOAD(conteiro);
				LCD_EN <= '1';
				LCD_RW <= '0';
				LCD_RS <= '1';
				
		WHEN LOAD_MSG_EN =>
				LCD_EN <= '0'; 
				LCD_RW <= '0';
				LCD_RS <= '1';
				
		WHEN LOAD_MENU_MSG =>
				LCD_DATA <= Linha_MSGOP_LOAD(conteiro);
				LCD_EN <= '1';
				LCD_RW <= '0';
				LCD_RS <= '1';
		
		WHEN LOAD_MENU_MSG_EN =>
				LCD_EN <= '0'; 
				LCD_RW <= '0';
				LCD_RS <= '1';

				
		WHEN NOT_MENU_MSG =>
				LCD_DATA <= Linha_MSGOP_NOT(conteiro);
				LCD_EN <= '1';
				LCD_RW <= '0';
				LCD_RS <= '1';
		
		WHEN NOT_MENU_MSG_EN =>
				LCD_EN <= '0'; 
				LCD_RW <= '0';
				LCD_RS <= '1';
				
		WHEN SWAP_MSG =>
				LCD_DATA <= Linha_SWAP(conteiro);
				LCD_EN <= '1';
				LCD_RW <= '0';
				LCD_RS <= '1';
				
		WHEN SWAP_MSG_EN =>
				LCD_EN <= '0'; 
				LCD_RW <= '0';
				LCD_RS <= '1';

		WHEN SWAP_MENU_MSG =>
				LCD_DATA <= Linha_MSGOP_SWAP(conteiro);
				LCD_EN <= '1';
				LCD_RW <= '0';
				LCD_RS <= '1';
		
		WHEN SWAP_MENU_MSG_EN =>
				LCD_EN <= '0'; 
				LCD_RW <= '0';
				LCD_RS <= '1';
				
		WHEN COMP_MENU_MSG =>
				LCD_DATA <= Linha_MSGOP_COMP(conteiro);
				LCD_EN <= '1';
				LCD_RW <= '0';
				LCD_RS <= '1';
		
		WHEN COMP_MENU_MSG_EN =>
				LCD_EN <= '0'; 
				LCD_RW <= '0';
				LCD_RS <= '1';
				
		WHEN SOMA_MSG =>
				LCD_DATA <= Linha_SOMA(conteiro);
				LCD_EN <= '1';
				LCD_RW <= '0';
				LCD_RS <= '1';
				
		WHEN SOMA_MSG_EN =>
				LCD_EN <= '0'; 
				LCD_RW <= '0';
				LCD_RS <= '1';
				
		WHEN SOMA_MENU_MSG =>
				LCD_DATA <= Linha_MSGOP_SOMA(conteiro);
				LCD_EN <= '1';
				LCD_RW <= '0';
				LCD_RS <= '1';
		
		WHEN SOMA_MENU_MSG_EN =>
				LCD_EN <= '0'; 
				LCD_RW <= '0';
				LCD_RS <= '1';
				
---------------------------------------------------------------
		WHEN WRITE_RXR1_SOMA=>
		LCD_DATA <= "11000101";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';
		
		WHEN WRITE_RXR1_ADDRESS1_SOMA=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';		
	
		WHEN WRITE_RXR1_1_SOMA=>
		LCD_DATA <= "00110001";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_RXR1_1_EN_SOMA=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';		
		
		WHEN WRITE_RXR1_ADDRESS2_SOMA=>
		LCD_DATA <= "11001000";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';		
		
		WHEN WRITE_RXR1_ADDRESS2_EN_SOMA=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';					
		
		WHEN WRITE_1_SOMA=>
		LCD_DATA <= "00110001";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_1_EN_SOMA=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';


		
		WHEN WRITE_RXR2_SOMA=>
		LCD_DATA <= "11000101";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';
		
		WHEN WRITE_RXR2_ADDRESS1_SOMA=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';		
	
		WHEN WRITE_RXR2_1_SOMA=>
		LCD_DATA <= "00110010";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_RXR2_1_EN_SOMA=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';		
		
		WHEN WRITE_RXR2_ADDRESS2_SOMA=>
		LCD_DATA <= "11001000";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';		
		
		WHEN WRITE_RXR2_ADDRESS2_EN_SOMA=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';					
		
		WHEN WRITE_2_SOMA=>
		LCD_DATA <= "00110010";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_2_EN_SOMA=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';

		
		
		WHEN WRITE_RXR3_SOMA=>
		LCD_DATA <= "11000101";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';
		
		WHEN WRITE_RXR3_ADDRESS1_SOMA=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';		
	
		WHEN WRITE_RXR3_1_SOMA=>
		LCD_DATA <= "00110011";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_RXR3_1_EN_SOMA=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';		
		
		WHEN WRITE_RXR3_ADDRESS2_SOMA=>
		LCD_DATA <= "11001000";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';		
		
		WHEN WRITE_RXR3_ADDRESS2_EN_SOMA=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';					
		
		WHEN WRITE_3_SOMA=>
		LCD_DATA <= "00110011";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_3_EN_SOMA=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		
		
		
		WHEN WRITE_RX_SOMA=>
		LCD_DATA <= "11000101";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';
		
		WHEN WRITE_RX_ADDRESS1_SOMA=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';		
	
		WHEN WRITE_RX_1_SOMA=>
		LCD_DATA <= "01111000";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_RX_1_EN_SOMA=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';		
		
		WHEN WRITE_RX_ADDRESS2_SOMA=>
		LCD_DATA <= "11001000";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';		
		
		WHEN WRITE_RX_ADDRESS2_EN_SOMA=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';					
		
		WHEN WRITE_x_SOMA=>
		LCD_DATA <= "01111000";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_x_EN_SOMA=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		
		
		WHEN WRITE_RYR1_SOMA=>
		LCD_DATA <= "11001011";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';
		
		WHEN WRITE_RYR1_ADDRESS1_SOMA=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';		
		
		WHEN WRITE_1Y_SOMA=>
		LCD_DATA <= "00110001";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_1Y_EN_SOMA =>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		
		WHEN WRITE_RYR2_SOMA=>
		LCD_DATA <= "11001011";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';
		
		WHEN WRITE_RYR2_ADDRESS1_SOMA=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';		
		
		WHEN WRITE_2Y_SOMA=>
		LCD_DATA <= "00110010";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_2Y_EN_SOMA =>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';

	
	
		WHEN WRITE_RYR3_SOMA=>
		LCD_DATA <= "11001011";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';
		
		WHEN WRITE_RYR3_ADDRESS1_SOMA=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';		
		
		WHEN WRITE_3Y_SOMA=>
		LCD_DATA <= "00110011";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_3Y_EN_SOMA =>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';

	
	
		WHEN WRITE_RY_SOMA=>
		LCD_DATA <= "11001011";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';
		
		WHEN WRITE_RY_ADDRESS1_SOMA=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';		
		
		WHEN WRITE_Y_SOMA=>
		LCD_DATA <= "01111001";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_Y_EN_SOMA =>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';
---------------------------------------------------------------
---------------------------------------------------------------
		WHEN WRITE_RXR1_SUB=>
		LCD_DATA <= "11000101";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';
		
		WHEN WRITE_RXR1_ADDRESS1_SUB=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';		
	
		WHEN WRITE_RXR1_1_SUB=>
		LCD_DATA <= "00110001";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_RXR1_1_EN_SUB=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';		
		
		WHEN WRITE_RXR1_ADDRESS2_SUB=>
		LCD_DATA <= "11001000";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';		
		
		WHEN WRITE_RXR1_ADDRESS2_EN_SUB=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';					
		
		WHEN WRITE_1_SUB=>
		LCD_DATA <= "00110001";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_1_EN_SUB=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';
	


		
		WHEN WRITE_RXR2_SUB=>
		LCD_DATA <= "11000101";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';
		
		WHEN WRITE_RXR2_ADDRESS1_SUB=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';		
	
		WHEN WRITE_RXR2_1_SUB=>
		LCD_DATA <= "00110010";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_RXR2_1_EN_SUB=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';		
		
		WHEN WRITE_RXR2_ADDRESS2_SUB=>
		LCD_DATA <= "11001000";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';		
		
		WHEN WRITE_RXR2_ADDRESS2_EN_SUB=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';					
		
		WHEN WRITE_2_SUB=>
		LCD_DATA <= "00110010";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_2_EN_SUB=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';

		
		
		WHEN WRITE_RXR3_SUB=>
		LCD_DATA <= "11000101";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';
		
		WHEN WRITE_RXR3_ADDRESS1_SUB=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';		
	
		WHEN WRITE_RXR3_1_SUB=>
		LCD_DATA <= "00110011";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_RXR3_1_EN_SUB=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';		
		
		WHEN WRITE_RXR3_ADDRESS2_SUB=>
		LCD_DATA <= "11001000";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';		
		
		WHEN WRITE_RXR3_ADDRESS2_EN_SUB=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';					
		
		WHEN WRITE_3_SUB=>
		LCD_DATA <= "00110011";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_3_EN_SUB=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		
		
		
		WHEN WRITE_RX_SUB=>
		LCD_DATA <= "11000101";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';
		
		WHEN WRITE_RX_ADDRESS1_SUB=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';		
	
		WHEN WRITE_RX_1_SUB=>
		LCD_DATA <= "01111000";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_RX_1_EN_SUB=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';		
		
		WHEN WRITE_RX_ADDRESS2_SUB=>
		LCD_DATA <= "11001000";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';		
		
		WHEN WRITE_RX_ADDRESS2_EN_SUB=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';					
		
		WHEN WRITE_x_SUB=>
		LCD_DATA <= "01111000";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_x_EN_SUB=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		
		
		WHEN WRITE_RYR1_SUB=>
		LCD_DATA <= "11001011";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';
		
		WHEN WRITE_RYR1_ADDRESS1_SUB=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';		
		
		WHEN WRITE_1Y_SUB=>
		LCD_DATA <= "00110001";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_1Y_EN_SUB =>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		
		WHEN WRITE_RYR2_SUB=>
		LCD_DATA <= "11001011";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';
		
		WHEN WRITE_RYR2_ADDRESS1_SUB=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';		
		
		WHEN WRITE_2Y_SUB=>
		LCD_DATA <= "00110010";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_2Y_EN_SUB =>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';

	
	
		WHEN WRITE_RYR3_SUB=>
		LCD_DATA <= "11001011";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';
		
		WHEN WRITE_RYR3_ADDRESS1_SUB=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';		
		
		WHEN WRITE_3Y_SUB=>
		LCD_DATA <= "00110011";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_3Y_EN_SUB =>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';

	
	
		WHEN WRITE_RY_SUB=>
		LCD_DATA <= "11001011";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';
		
		WHEN WRITE_RY_ADDRESS1_SUB=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';		
		
		WHEN WRITE_Y_SUB=>
		LCD_DATA <= "01111001";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_Y_EN_SUB =>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';
---------------------------------------------------------------
---------------------------------------------------------------
		WHEN WRITE_RXR1_AND=>
		LCD_DATA <= "11000101";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';
		
		WHEN WRITE_RXR1_ADDRESS1_AND=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';		
	
		WHEN WRITE_RXR1_1_AND=>
		LCD_DATA <= "00110001";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_RXR1_1_EN_AND=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';		
		
		WHEN WRITE_RXR1_ADDRESS2_AND=>
		LCD_DATA <= "11001000";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';		
		
		WHEN WRITE_RXR1_ADDRESS2_EN_AND=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';					
		
		WHEN WRITE_1_AND=>
		LCD_DATA <= "00110001";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_1_EN_AND=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';


		
		WHEN WRITE_RXR2_AND=>
		LCD_DATA <= "11000101";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';
		
		WHEN WRITE_RXR2_ADDRESS1_AND=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';		
	
		WHEN WRITE_RXR2_1_AND=>
		LCD_DATA <= "00110010";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_RXR2_1_EN_AND=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';		
		
		WHEN WRITE_RXR2_ADDRESS2_AND=>
		LCD_DATA <= "11001000";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';		
		
		WHEN WRITE_RXR2_ADDRESS2_EN_AND=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';					
		
		WHEN WRITE_2_AND=>
		LCD_DATA <= "00110010";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_2_EN_AND=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';

		
		
		WHEN WRITE_RXR3_AND=>
		LCD_DATA <= "11000101";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';
		
		WHEN WRITE_RXR3_ADDRESS1_AND=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';		
	
		WHEN WRITE_RXR3_1_AND=>
		LCD_DATA <= "00110011";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_RXR3_1_EN_AND=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';		
		
		WHEN WRITE_RXR3_ADDRESS2_AND=>
		LCD_DATA <= "11001000";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';		
		
		WHEN WRITE_RXR3_ADDRESS2_EN_AND=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';					
		
		WHEN WRITE_3_AND=>
		LCD_DATA <= "00110011";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_3_EN_AND=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		
		
		
		WHEN WRITE_RX_AND=>
		LCD_DATA <= "11000101";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';
		
		WHEN WRITE_RX_ADDRESS1_AND=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';		
	
		WHEN WRITE_RX_1_AND=>
		LCD_DATA <= "01111000";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_RX_1_EN_AND=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';		
		
		WHEN WRITE_RX_ADDRESS2_AND=>
		LCD_DATA <= "11001000";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';		
		
		WHEN WRITE_RX_ADDRESS2_EN_AND=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';					
		
		WHEN WRITE_x_AND=>
		LCD_DATA <= "01111000";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_x_EN_AND=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		
		
		WHEN WRITE_RYR1_AND=>
		LCD_DATA <= "11001011";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';
		
		WHEN WRITE_RYR1_ADDRESS1_AND=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';		
		
		WHEN WRITE_1Y_AND=>
		LCD_DATA <= "00110001";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_1Y_EN_AND =>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		
		WHEN WRITE_RYR2_AND=>
		LCD_DATA <= "11001011";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';
		
		WHEN WRITE_RYR2_ADDRESS1_AND=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';		
		
		WHEN WRITE_2Y_AND=>
		LCD_DATA <= "00110010";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_2Y_EN_AND =>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';

	
	
		WHEN WRITE_RYR3_AND=>
		LCD_DATA <= "11001011";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';
		
		WHEN WRITE_RYR3_ADDRESS1_AND=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';		
		
		WHEN WRITE_3Y_AND=>
		LCD_DATA <= "00110011";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_3Y_EN_AND =>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';

	
	
		WHEN WRITE_RY_AND=>
		LCD_DATA <= "11001011";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';
		
		WHEN WRITE_RY_ADDRESS1_AND=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';		
		
		WHEN WRITE_Y_AND=>
		LCD_DATA <= "01111001";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_Y_EN_AND =>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';
---------------------------------------------------------------
---------------------------------------------------------------
		WHEN WRITE_RXR1_OR=>
		LCD_DATA <= "11000101";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';
		
		WHEN WRITE_RXR1_ADDRESS1_OR=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';		
	
		WHEN WRITE_RXR1_1_OR=>
		LCD_DATA <= "00110001";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_RXR1_1_EN_OR=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';		
		
		WHEN WRITE_RXR1_ADDRESS2_OR=>
		LCD_DATA <= "11001000";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';		
		
		WHEN WRITE_RXR1_ADDRESS2_EN_OR=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';					
		
		WHEN WRITE_1_OR=>
		LCD_DATA <= "00110001";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_1_EN_OR=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';


		
		WHEN WRITE_RXR2_OR=>
		LCD_DATA <= "11000101";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';
		
		WHEN WRITE_RXR2_ADDRESS1_OR=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';		
	
		WHEN WRITE_RXR2_1_OR=>
		LCD_DATA <= "00110010";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_RXR2_1_EN_OR=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';		
		
		WHEN WRITE_RXR2_ADDRESS2_OR=>
		LCD_DATA <= "11001000";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';		
		
		WHEN WRITE_RXR2_ADDRESS2_EN_OR=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';					
		
		WHEN WRITE_2_OR=>
		LCD_DATA <= "00110010";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_2_EN_OR=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';

		
		
		WHEN WRITE_RXR3_OR=>
		LCD_DATA <= "11000101";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';
		
		WHEN WRITE_RXR3_ADDRESS1_OR=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';		
	
		WHEN WRITE_RXR3_1_OR=>
		LCD_DATA <= "00110011";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_RXR3_1_EN_OR=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';		
		
		WHEN WRITE_RXR3_ADDRESS2_OR=>
		LCD_DATA <= "11001000";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';		
		
		WHEN WRITE_RXR3_ADDRESS2_EN_OR=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';					
		
		WHEN WRITE_3_OR=>
		LCD_DATA <= "00110011";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_3_EN_OR=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		
		
		
		WHEN WRITE_RX_OR=>
		LCD_DATA <= "11000101";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';
		
		WHEN WRITE_RX_ADDRESS1_OR=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';		
	
		WHEN WRITE_RX_1_OR=>
		LCD_DATA <= "01111000";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_RX_1_EN_OR=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';		
		
		WHEN WRITE_RX_ADDRESS2_OR=>
		LCD_DATA <= "11001000";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';		
		
		WHEN WRITE_RX_ADDRESS2_EN_OR=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';					
		
		WHEN WRITE_x_OR=>
		LCD_DATA <= "01111000";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_x_EN_OR=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		
		
		WHEN WRITE_RYR1_OR=>
		LCD_DATA <= "11001011";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';
		
		WHEN WRITE_RYR1_ADDRESS1_OR=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';		
		
		WHEN WRITE_1Y_OR=>
		LCD_DATA <= "00110001";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_1Y_EN_OR =>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		
		WHEN WRITE_RYR2_OR=>
		LCD_DATA <= "11001011";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';
		
		WHEN WRITE_RYR2_ADDRESS1_OR=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';		
		
		WHEN WRITE_2Y_OR=>
		LCD_DATA <= "00110010";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_2Y_EN_OR =>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';

	
	
		WHEN WRITE_RYR3_OR=>
		LCD_DATA <= "11001011";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';
		
		WHEN WRITE_RYR3_ADDRESS1_OR=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';		
		
		WHEN WRITE_3Y_OR=>
		LCD_DATA <= "00110011";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_3Y_EN_OR =>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';

	
	
		WHEN WRITE_RY_OR=>
		LCD_DATA <= "11001011";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';
		
		WHEN WRITE_RY_ADDRESS1_OR=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';		
		
		WHEN WRITE_Y_OR=>
		LCD_DATA <= "01111001";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_Y_EN_OR =>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';
---------------------------------------------------------------
---------------------------------------------------------------
		WHEN WRITE_RXR1_MUL=>
		LCD_DATA <= "11000101";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';
		
		WHEN WRITE_RXR1_ADDRESS1_MUL=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';		
	
		WHEN WRITE_RXR1_1_MUL=>
		LCD_DATA <= "00110001";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_RXR1_1_EN_MUL=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';		
		
		WHEN WRITE_RXR1_ADDRESS2_MUL=>
		LCD_DATA <= "11001000";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';		
		
		WHEN WRITE_RXR1_ADDRESS2_EN_MUL=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';					
		
		WHEN WRITE_1_MUL=>
		LCD_DATA <= "00110001";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_1_EN_MUL=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';
	


		
		WHEN WRITE_RXR2_MUL=>
		LCD_DATA <= "11000101";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';
		
		WHEN WRITE_RXR2_ADDRESS1_MUL=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';		
	
		WHEN WRITE_RXR2_1_MUL=>
		LCD_DATA <= "00110010";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_RXR2_1_EN_MUL=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';		
		
		WHEN WRITE_RXR2_ADDRESS2_MUL=>
		LCD_DATA <= "11001000";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';		
		
		WHEN WRITE_RXR2_ADDRESS2_EN_MUL=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';					
		
		WHEN WRITE_2_MUL=>
		LCD_DATA <= "00110010";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_2_EN_MUL=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';

		
		
		WHEN WRITE_RXR3_MUL=>
		LCD_DATA <= "11000101";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';
		
		WHEN WRITE_RXR3_ADDRESS1_MUL=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';		
	
		WHEN WRITE_RXR3_1_MUL=>
		LCD_DATA <= "00110011";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_RXR3_1_EN_MUL=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';		
		
		WHEN WRITE_RXR3_ADDRESS2_MUL=>
		LCD_DATA <= "11001000";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';		
		
		WHEN WRITE_RXR3_ADDRESS2_EN_MUL=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';					
		
		WHEN WRITE_3_MUL=>
		LCD_DATA <= "00110011";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_3_EN_MUL=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		
		
		
		WHEN WRITE_RX_MUL=>
		LCD_DATA <= "11000101";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';
		
		WHEN WRITE_RX_ADDRESS1_MUL=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';		
	
		WHEN WRITE_RX_1_MUL=>
		LCD_DATA <= "01111000";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_RX_1_EN_MUL=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';		
		
		WHEN WRITE_RX_ADDRESS2_MUL=>
		LCD_DATA <= "11001000";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';		
		
		WHEN WRITE_RX_ADDRESS2_EN_MUL=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';					
		
		WHEN WRITE_x_MUL=>
		LCD_DATA <= "01111000";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_x_EN_MUL=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		
		
		WHEN WRITE_RYR1_MUL=>
		LCD_DATA <= "11001011";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';
		
		WHEN WRITE_RYR1_ADDRESS1_MUL=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';		
		
		WHEN WRITE_1Y_MUL=>
		LCD_DATA <= "00110001";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_1Y_EN_MUL =>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		
		WHEN WRITE_RYR2_MUL=>
		LCD_DATA <= "11001011";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';
		
		WHEN WRITE_RYR2_ADDRESS1_MUL=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';		
		
		WHEN WRITE_2Y_MUL=>
		LCD_DATA <= "00110010";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_2Y_EN_MUL =>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';

	
	
		WHEN WRITE_RYR3_MUL=>
		LCD_DATA <= "11001011";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';
		
		WHEN WRITE_RYR3_ADDRESS1_MUL=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';		
		
		WHEN WRITE_3Y_MUL=>
		LCD_DATA <= "00110011";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_3Y_EN_MUL =>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';

	
	
		WHEN WRITE_RY_MUL=>
		LCD_DATA <= "11001011";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';
		
		WHEN WRITE_RY_ADDRESS1_MUL=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';		
		
		WHEN WRITE_Y_MUL=>
		LCD_DATA <= "01111001";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_Y_EN_MUL =>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';
---------------------------------------------------------------
---------------------------------------------------------------
		WHEN WRITE_RYR1_LOAD=>
		LCD_DATA <= "11000101";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';
		
		WHEN WRITE_RYR1_ADDRESS1_LOAD=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';		
		
		WHEN WRITE_1Y_LOAD=>
		LCD_DATA <= "00110001";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_1Y_EN_LOAD =>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		
		WHEN WRITE_RYR2_LOAD=>
		LCD_DATA <= "11000101";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';
		
		WHEN WRITE_RYR2_ADDRESS1_LOAD=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';		
		
		WHEN WRITE_2Y_LOAD=>
		LCD_DATA <= "00110010";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_2Y_EN_LOAD =>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';

	
	
		WHEN WRITE_RYR3_LOAD=>
		LCD_DATA <= "11000101";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';
		
		WHEN WRITE_RYR3_ADDRESS1_LOAD=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';		
		
		WHEN WRITE_3Y_LOAD=>
		LCD_DATA <= "00110011";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_3Y_EN_LOAD =>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';

	
	
		WHEN WRITE_RY_LOAD=>
		LCD_DATA <= "11000101";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';
		
		WHEN WRITE_RY_ADDRESS1_LOAD=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';		
		
		WHEN WRITE_Y_LOAD=>
		LCD_DATA <= "01111001";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_Y_EN_LOAD =>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';
---------------------------------------------------------------
---------------------------------------------------------------
		WHEN WRITE_RXR1_NOT=>
		LCD_DATA <= "11000110";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';
		
		WHEN WRITE_RXR1_ADDRESS1_NOT=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';		
		
		WHEN WRITE_RXR1_1_NOT=>
		LCD_DATA <= "00110001";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_RXR1_1_EN_NOT =>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		
		WHEN WRITE_RXR2_NOT=>
		LCD_DATA <= "11000110";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';
		
		WHEN WRITE_RXR2_ADDRESS1_NOT=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';		
		
		WHEN WRITE_RXR2_1_NOT=>
		LCD_DATA <= "00110010";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_RXR2_1_EN_NOT=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';

	
	
		WHEN WRITE_RXR3_NOT=>
		LCD_DATA <= "11000110";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';
		
		WHEN WRITE_RXR3_ADDRESS1_NOT=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';		
		
		WHEN WRITE_RXR3_1_NOT=>
		LCD_DATA <= "00110011";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_RXR3_1_EN_NOT =>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';

	
	
		WHEN WRITE_RX_NOT=>
		LCD_DATA <= "11000110";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';
		
		WHEN WRITE_RX_ADDRESS1_NOT=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';		
		
		WHEN WRITE_RX_1_NOT=>
		LCD_DATA <= "01111000";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_RX_1_EN_NOT=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';



		WHEN WRITE_RYR1_NOT=>
		LCD_DATA <= "11001010";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';
		
		WHEN WRITE_RYR1_ADDRESS1_NOT=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';		
		
		WHEN WRITE_RYR1_1_NOT=>
		LCD_DATA <= "00110001";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_RYR1_1_EN_NOT =>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		
		WHEN WRITE_RYR2_NOT=>
		LCD_DATA <= "11001010";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';
		
		WHEN WRITE_RYR2_ADDRESS1_NOT=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';		
		
		WHEN WRITE_RYR2_1_NOT=>
		LCD_DATA <= "00110010";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_RYR2_1_EN_NOT=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';

	
	
		WHEN WRITE_RYR3_NOT=>
		LCD_DATA <= "11001010";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';
		
		WHEN WRITE_RYR3_ADDRESS1_NOT=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';		
		
		WHEN WRITE_RYR3_1_NOT=>
		LCD_DATA <= "00110011";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_RYR3_1_EN_NOT =>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';

	
	
		WHEN WRITE_RY_NOT=>
		LCD_DATA <= "11001010";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';
		
		WHEN WRITE_RY_ADDRESS1_NOT=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';		
		
		WHEN WRITE_RY_1_NOT=>
		LCD_DATA <= "01111001";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_RY_1_EN_NOT=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';
---------------------------------------------------------------
---------------------------------------------------------------
		WHEN WRITE_RXR1_SWAP=>
		LCD_DATA <= "11000110";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';
		
		WHEN WRITE_RXR1_ADDRESS1_SWAP=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';		
		
		WHEN WRITE_RXR1_1_SWAP=>
		LCD_DATA <= "00110001";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_RXR1_1_EN_SWAP=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		
		WHEN WRITE_RXR2_SWAP=>
		LCD_DATA <= "11000110";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';
		
		WHEN WRITE_RXR2_ADDRESS1_SWAP=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';		
		
		WHEN WRITE_RXR2_1_SWAP=>
		LCD_DATA <= "00110010";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_RXR2_1_EN_SWAP=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';

	
	
		WHEN WRITE_RXR3_SWAP=>
		LCD_DATA <= "11000110";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';
		
		WHEN WRITE_RXR3_ADDRESS1_SWAP=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';		
		
		WHEN WRITE_RXR3_1_SWAP=>
		LCD_DATA <= "00110011";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_RXR3_1_EN_SWAP=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';

	
	
		WHEN WRITE_RX_SWAP=>
		LCD_DATA <= "11000110";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';
		
		WHEN WRITE_RX_ADDRESS1_SWAP=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';		
		
		WHEN WRITE_RX_1_SWAP=>
		LCD_DATA <= "01111000";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_RX_1_EN_SWAP=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';



		WHEN WRITE_RYR1_SWAP=>
		LCD_DATA <= "11001010";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';
		
		WHEN WRITE_RYR1_ADDRESS1_SWAP=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';		
		
		WHEN WRITE_RYR1_1_SWAP=>
		LCD_DATA <= "00110001";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_RYR1_1_EN_SWAP=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		
		WHEN WRITE_RYR2_SWAP=>
		LCD_DATA <= "11001010";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';
		
		WHEN WRITE_RYR2_ADDRESS1_SWAP=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';		
		
		WHEN WRITE_RYR2_1_SWAP=>
		LCD_DATA <= "00110010";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_RYR2_1_EN_SWAP=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';

	
	
		WHEN WRITE_RYR3_SWAP=>
		LCD_DATA <= "11001010";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';
		
		WHEN WRITE_RYR3_ADDRESS1_SWAP=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';		
		
		WHEN WRITE_RYR3_1_SWAP=>
		LCD_DATA <= "00110011";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_RYR3_1_EN_SWAP=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';

	
	
		WHEN WRITE_RY_SWAP=>
		LCD_DATA <= "11001010";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';
		
		WHEN WRITE_RY_ADDRESS1_SWAP=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';		
		
		WHEN WRITE_RY_1_SWAP=>
		LCD_DATA <= "01111001";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_RY_1_EN_SWAP=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';
---------------------------------------------------------------
---------------------------------------------------------------
---------------------------------------------------------------
		WHEN WRITE_RXR1_COMP=>
		LCD_DATA <= "11000110";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';
		
		WHEN WRITE_RXR1_ADDRESS1_COMP=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';		
		
		WHEN WRITE_RXR1_1_COMP=>
		LCD_DATA <= "00110001";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_RXR1_1_EN_COMP=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		
		WHEN WRITE_RXR2_COMP=>
		LCD_DATA <= "11000110";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';
		
		WHEN WRITE_RXR2_ADDRESS1_COMP=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';		
		
		WHEN WRITE_RXR2_1_COMP=>
		LCD_DATA <= "00110010";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_RXR2_1_EN_COMP=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';

	
	
		WHEN WRITE_RXR3_COMP=>
		LCD_DATA <= "11000110";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';
		
		WHEN WRITE_RXR3_ADDRESS1_COMP=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';		
		
		WHEN WRITE_RXR3_1_COMP=>
		LCD_DATA <= "00110011";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_RXR3_1_EN_COMP=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';

	
	
		WHEN WRITE_RX_COMP=>
		LCD_DATA <= "11000110";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';
		
		WHEN WRITE_RX_ADDRESS1_COMP=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';		
		
		WHEN WRITE_RX_1_COMP=>
		LCD_DATA <= "01111000";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_RX_1_EN_COMP=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';



		WHEN WRITE_RYR1_COMP=>
		LCD_DATA <= "11001001";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';
		
		WHEN WRITE_RYR1_ADDRESS1_COMP=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';		
		
		WHEN WRITE_RYR1_1_COMP=>
		LCD_DATA <= "00110001";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_RYR1_1_EN_COMP=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		
		WHEN WRITE_RYR2_COMP=>
		LCD_DATA <= "11001001";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';
		
		WHEN WRITE_RYR2_ADDRESS1_COMP=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';		
		
		WHEN WRITE_RYR2_1_COMP=>
		LCD_DATA <= "00110010";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_RYR2_1_EN_COMP=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';

	
	
		WHEN WRITE_RYR3_COMP=>
		LCD_DATA <= "11001001";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';
		
		WHEN WRITE_RYR3_ADDRESS1_COMP=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';		
		
		WHEN WRITE_RYR3_1_COMP=>
		LCD_DATA <= "00110011";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_RYR3_1_EN_COMP=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';

	
	
		WHEN WRITE_RY_COMP=>
		LCD_DATA <= "11001001";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';
		
		WHEN WRITE_RY_ADDRESS1_COMP=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';		
		
		WHEN WRITE_RY_1_COMP=>
		LCD_DATA <= "01111001";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN WRITE_RY_1_EN_COMP=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		
		
		WHEN COMP_ADDRESS_OPERATOR=>
		LCD_DATA <= "11000111";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '0';
		
		WHEN COMP_ADDRESS_OPERATOR_EN=>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '0';	
		
		
		WHEN COMP_WAIT =>
		LCD_DATA <= "00111111";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN COMP_WAIT_EN =>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		
		WHEN COMP_MAIOR =>
		LCD_DATA <= "00111110";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';	
	
		WHEN COMP_MAIOR_EN =>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		
		WHEN COMP_MENOR =>
		LCD_DATA <= "00111100";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';	
		
		WHEN COMP_MENOR_EN =>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';
		
		WHEN COMP_IGUAL =>
		LCD_DATA <= "00111101";
		LCD_EN <= '1';
		LCD_RW <= '0';
		LCD_RS <= '1';	
		
		WHEN COMP_IGUAL_EN =>
		LCD_EN <= '0';
		LCD_RW <= '0';
		LCD_RS <= '1';
---------------------------------------------------------------
		WHEN SUB_MSG =>
				LCD_DATA <= Linha_SUB(conteiro);
				LCD_EN <= '1';
				LCD_RW <= '0';
				LCD_RS <= '1';
				
		WHEN SUB_MSG_EN =>
				LCD_EN <= '0'; 
				LCD_RW <= '0';
				LCD_RS <= '1';
				
		WHEN SUB_MENU_MSG =>
				LCD_DATA <= Linha_MSGOP_SUB(conteiro);
				LCD_EN <= '1';
				LCD_RW <= '0';
				LCD_RS <= '1';
		
		WHEN SUB_MENU_MSG_EN =>
				LCD_EN <= '0'; 
				LCD_RW <= '0';
				LCD_RS <= '1';
				
				
		WHEN AND_MSG =>
				LCD_DATA <= Linha_AND(conteiro);
				LCD_EN <= '1';
				LCD_RW <= '0';
				LCD_RS <= '1';
				
		WHEN AND_MSG_EN =>
				LCD_EN <= '0'; 
				LCD_RW <= '0';
				LCD_RS <= '1';

		WHEN AND_MENU_MSG =>
				LCD_DATA <= Linha_MSGOP_AND(conteiro);
				LCD_EN <= '1';
				LCD_RW <= '0';
				LCD_RS <= '1';
		
		WHEN AND_MENU_MSG_EN =>
				LCD_EN <= '0'; 
				LCD_RW <= '0';
				LCD_RS <= '1';

				
		WHEN NOT_MSG =>
				LCD_DATA <= Linha_NOT(conteiro);
				LCD_EN <= '1';
				LCD_RW <= '0';
				LCD_RS <= '1';
				
		WHEN NOT_MSG_EN =>
				LCD_EN <= '0'; 
				LCD_RW <= '0';
				LCD_RS <= '1';

				
		WHEN OR_MSG =>
				LCD_DATA <= Linha_OR(conteiro);
				LCD_EN <= '1';
				LCD_RW <= '0';
				LCD_RS <= '1';
				
		WHEN OR_MSG_EN =>
				LCD_EN <= '0'; 
				LCD_RW <= '0';
				LCD_RS <= '1';

		WHEN OR_MENU_MSG =>
				LCD_DATA <= Linha_MSGOP_OR(conteiro);
				LCD_EN <= '1';
				LCD_RW <= '0';
				LCD_RS <= '1';
		
		WHEN OR_MENU_MSG_EN =>
				LCD_EN <= '0'; 
				LCD_RW <= '0';
				LCD_RS <= '1';

		WHEN COMP_MSG =>
				LCD_DATA <= Linha_COMP(conteiro);
				LCD_EN <= '1';
				LCD_RW <= '0';
				LCD_RS <= '1';
				
		WHEN COMP_MSG_EN =>
				LCD_EN <= '0'; 
				LCD_RW <= '0';
				LCD_RS <= '1';

				
		WHEN MUL_MSG =>
				LCD_DATA <= Linha_MULT(conteiro);
				LCD_EN <= '1';
				LCD_RW <= '0';
				LCD_RS <= '1';
				
		WHEN MUL_MSG_EN =>
				LCD_EN <= '0'; 
				LCD_RW <= '0';
				LCD_RS <= '1';
				
				
		WHEN MUL_MENU_MSG =>
				LCD_DATA <= Linha_MSGOP_MUL(conteiro);
				LCD_EN <= '1';
				LCD_RW <= '0';
				LCD_RS <= '1';
		
		WHEN MUL_MENU_MSG_EN =>
				LCD_EN <= '0'; 
				LCD_RW <= '0';
				LCD_RS <= '1';
				
		WHEN MENU_MSG =>
				LCD_DATA <= Linha_MENU(conteiro);
				LCD_EN <= '1';
				LCD_RW <= '0';
				LCD_RS <= '1';
				
		WHEN MENU_MSG_EN =>
				LCD_EN <= '0'; 
				LCD_RW <= '0';
				LCD_RS <= '1';
		WHEN OTHERS =>
			NULL;

			END CASE;
END PROCESS;



END bhv;