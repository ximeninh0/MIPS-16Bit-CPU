LIBRARY ieee;
USE ieee.std_logic_1164.all;
use work.CPU_PACKAGE.all;

ENTITY PIPE_ID_EX IS 
    port(
        -- Inputs
        A_IN : IN STD_LOGIC_VECTOR(15 DOWNTO 0); -- Registrador A (rs)
        B_IN : IN STD_LOGIC_VECTOR(15 DOWNTO 0); -- Registrador B (rt)
        SIGNAL_EXT_IN : IN STD_LOGIC_VECTOR(15 DOWNTO 0); -- Imediato estendido
        IF_ID_REG_RS_IN : IN STD_LOGIC_VECTOR(3 DOWNTO 0); -- Código do registrador rs
        IF_ID_REG_RT_IN : IN STD_LOGIC_VECTOR(3 DOWNTO 0); -- Código do registrador rt
        IF_ID_REG_RD_IN : IN STD_LOGIC_VECTOR(3 DOWNTO 0); -- Código do registrador rd
        NEXT_PC_IN : IN STD_LOGIC_VECTOR(15 DOWNTO 0); -- Próximo PC

        -- Outputs
        A_OUT : OUT STD_LOGIC_VECTOR(15 DOWNTO 0); -- Registrador A (rs)
        B_OUT : OUT STD_LOGIC_VECTOR(15 DOWNTO 0); -- Registrador B (rt)
        SIGNAL_EXT_OUT : OUT STD_LOGIC_VECTOR(15 DOWNTO 0); -- Imediato estendido
        IF_ID_REG_RS_OUT : OUT STD_LOGIC_VECTOR(3 DOWNTO 0); -- Código do registrador rs
        IF_ID_REG_RT_OUT : OUT STD_LOGIC_VECTOR(3 DOWNTO 0); -- Código do registrador rt
        IF_ID_REG_RD_OUT : OUT STD_LOGIC_VECTOR(3 DOWNTO 0); -- Código do registrador rd
        NEXT_PC_OUT : OUT STD_LOGIC_VECTOR(15 DOWNTO 0); -- Próximo PC

        -- Sinais de controle
        -- EX
        EX_ALU_SRC_IN : IN STD_LOGIC;
        EX_REG_DST_IN : IN STD_LOGIC;
        EX_ALU_OP_IN : IN STD_LOGIC_VECTOR(1 DOWNTO 0);

        EX_ALU_SRC_OUT : OUT STD_LOGIC;
        EX_REG_DST_OUT : OUT STD_LOGIC;
        EX_ALU_OP_OUT : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);

        -- MEM
        MEM_WRITE_IN : IN STD_LOGIC;
        MEM_READ_IN : IN STD_LOGIC;
        -- MEM_ALU_RESULT_IN : IN STD_LOGIC;
        -- MEM_ALU_SRC2_IN : IN STD_LOGIC;

        MEM_WRITE_OUT : OUT STD_LOGIC;
        MEM_READ_OUT : OUT STD_LOGIC;
        -- MEM_ALU_RESULT_OUT : OUT STD_LOGIC;
        -- MEM_ALU_SRC2_OUT : OUT STD_LOGIC;

        -- WB
        WB_MEM_TO_REG_IN : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
        WB_REG_WRITE_IN : IN STD_LOGIC;

        WB_MEM_TO_REG_OUT : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
        WB_REG_WRITE_OUT : OUT STD_LOGIC;

        -- Controle de clock e reset
        CLOCK : IN STD_LOGIC;
        RESET : IN STD_LOGIC

    );
END PIPE_ID_EX;


ARCHITECTURE Behavior OF PIPE_ID_EX IS
	BEGIN
    -- Instanciação dos registradores do estágio ID/EX
    REG_A_INSTANCE: LOW_WRITE_REG16 PORT MAP(A_IN,'1',RESET,CLOCK,A_OUT);
	 REG_B_INSTANCE: LOW_WRITE_REG16 PORT MAP(B_IN,'1',RESET,CLOCK,B_OUT);
    SIGNAL_EXT_INSTANCE: LOW_WRITE_REG16 PORT MAP(SIGNAL_EXT_IN,'1',RESET,CLOCK,SIGNAL_EXT_OUT);

    IF_ID_REG_RS_INSTANCE: FOUR_BIT_REG PORT MAP(IF_ID_REG_RS_IN,'1',RESET,CLOCK,IF_ID_REG_RS_OUT);
    IF_ID_REG_RT_INSTANCE: FOUR_BIT_REG PORT MAP(IF_ID_REG_RT_IN,'1',RESET,CLOCK,IF_ID_REG_RT_OUT);
	 IF_ID_REG_RD_INSTANCE: FOUR_BIT_REG PORT MAP(IF_ID_REG_RD_IN,'1',RESET,CLOCK,IF_ID_REG_RD_OUT);


    NEXT_PC_INSTANCE: REG PORT MAP(NEXT_PC_IN,'1',RESET,CLOCK,NEXT_PC_OUT);

    -- Sinais de controle
    -- EX
    EX_ALU_SRC_INSTANCE: ONE_BIT_REG PORT MAP(EX_ALU_SRC_IN,'1',RESET,CLOCK,EX_ALU_SRC_OUT);
    EX_REG_DST_INSTANCE: ONE_BIT_REG PORT MAP(EX_REG_DST_IN,'1',RESET,CLOCK,EX_REG_DST_OUT);
    EX_ALU_OP_INSTANCE: TWO_BIT_REG PORT MAP(EX_ALU_OP_IN,'1',RESET,CLOCK,EX_ALU_OP_OUT);

    -- MEM
    MEM_WRITE_INSTANCE: ONE_BIT_REG PORT MAP(MEM_WRITE_IN,'1',RESET,CLOCK,MEM_WRITE_OUT);
    MEM_READ_INSTANCE: ONE_BIT_REG PORT MAP(MEM_READ_IN,'1',RESET,CLOCK,MEM_READ_OUT);
    -- MEM_ALU_RESULT_INSTANCE: ONE_BIT_REG PORT MAP(MEM_ALU_RESULT_IN,'1',RESET,CLOCK,MEM_ALU_RESULT_OUT);
    -- MEM_ALU_SRC2_INSTANCE: ONE_BIT_REG PORT MAP(MEM_ALU_SRC2_IN,'1',RESET,CLOCK,MEM_ALU_SRC2_OUT);

    -- WB
    WB_MEM_TO_REG_INSTANCE: TWO_BIT_REG PORT MAP(WB_MEM_TO_REG_IN,'1',RESET,CLOCK,WB_MEM_TO_REG_OUT);
    WB_REG_WRITE_INSTANCE: ONE_BIT_REG PORT MAP(WB_REG_WRITE_IN,'1',RESET,CLOCK,WB_REG_WRITE_OUT);


END Behavior;
