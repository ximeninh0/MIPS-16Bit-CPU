LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY AND_COMPONENT IS 
port(
	X,Y :IN std_logic_vector(3 DOWNTO 0);
	Z : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END AND_COMPONENT;

ARCHITECTURE Behavior OF AND_COMPONENT IS
-- SAIDA RECEBE AND ENTRE AS DUAS PORTAS
BEGIN
	Z <= X AND Y;

END Behavior;
