LIBRARY ieee;
USE ieee.std_logic_1164.all;
use work.CPU_PACKAGE.all;

ENTITY CPU IS 
	port(
		SW : IN STD_LOGIC_VECTOR(17 DOWNTO 0); -- Sinais de entrada e CLOCK da placa
		KEY: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		Clock_50 : IN STD_LOGIC;
		
		HEX0,HEX1,HEX2 : OUT STD_LOGIC_VECTOR(0 TO 6); -- Sinais de saída para os displays de 7 segmentos
		HEX4 : OUT STD_LOGIC_VECTOR(0 TO 6);
		HEX7 : OUT STD_LOGIC_VECTOR(0 TO 6);
		
		LEDR : OUT STD_LOGIC_VECTOR(17 DOWNTO 0);		-- Sinais de saída para os LEDS da placa
		LEDG: OUT STD_LOGIC_VECTOR(8 DOWNTO 0);
		
		LCD_DATA : out STD_LOGIC_VECTOR(7 DOWNTO 0); -- Sinais para manipulação do display LCD da placa
		LCD_RW : OUT STD_LOGIC;
		LCD_EN : OUT STD_LOGIC;
		LCD_RS: OUT STD_LOGIC
	);
END CPU;

ARCHITECTURE Behavior OF CPU IS

CONSTANT max: INTEGER := 500000;				-- Ciclo do clock (é ajustável)
CONSTANT half: INTEGER := max/2;				-- Meio Ciclo
SIGNAL clockticks: INTEGER RANGE 0 TO max;-- Conta cada ciclo do clock de entrada
SIGNAL CLOCK: STD_LOGIC;						-- Clock instanciado

SIGNAL RESET: STD_LOGIC := '0';				-- Sinal de reset geral

-- Sinais do Estagio IF
SIGNAL IF_PC_NEXT,IF_PC_CURRENT, IF_PC_MUX,IF_INSTRUCTION : STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL IF_PC_ADD_OVERFLOW, IF_PC_ADD_COUT : STD_LOGIC;
SIGNAL IF_NEXT_PC : STD_LOGIC_VECTOR(15 DOWNTO 0);

-- Sinais do Estagio IF/ID
SIGNAL ID_PC_SOURCE : STD_LOGIC_VECTOR(1 DOWNTO 0);
SIGNAL ID_IF_ID_WRITE, ID_PC_WRITE : STD_LOGIC;
SIGNAL ID_IF_FLUSH : STD_LOGIC;
SIGNAL ID_NEXT_PC : STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL ID_INSTRUCTION_DATA : STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL ID_SIGNAL_EXTENDED, ID_SIGNAL_SHIFTED : STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL ID_RS_OP, ID_RT_OP, ID_RD_OP : STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL ID_REG_DATA1, ID_REG_DATA2 : STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL ID_REG_EQUAL : STD_LOGIC;
SIGNAL ID_JUMP_ADDRESS : STD_LOGIC_VECTOR(15 DOWNTO 0); 
SIGNAL ID_RIPPLE_BRANCH_OVERFLOW, ID_RIPPLE_BRANCH_COUT : STD_LOGIC;
SIGNAL ID_BRANCH_RESULT : STD_LOGIC_VECTOR(15 DOWNTO 0);

SIGNAL ID_ALU_SRC, ID_REG_DST : STD_LOGIC;
SIGNAL ID_ALU_OP : STD_LOGIC_VECTOR(2 DOWNTO 0);
SIGNAL ID_MEM_WRITE, ID_MEM_READ, ID_MEM_TO_REG, ID_REG_WRITE : STD_LOGIC;
SIGNAL ID_IF_FLUSH, ID_ID_FLUSH, ID_EX_FLUSH, ID_WB_FLUSH : STD_LOGIC;

-- Sinais do Estagio ID/EX
SIGNAL EX_A, EX_B : STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL EX_SIGNAL_EXTENDED : STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL EX_RS_OP, EX_RT_OP, EX_RD_OP : STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL EX_NEXT_PC : STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL EX_ALU_SRC, EX_REG_DST : STD_LOGIC;
SIGNAL EX_ALU_OP : STD_LOGIC_VECTOR(1 DOWNTO 0);
SIGNAL EX_MEM_WRITE, EX_MEM_READ : STD_LOGIC;
SIGNAL EX_REG_WRITE : STD_LOGIC;
SIGNAL EX_MEM_TO_REG : STD_LOGIC_VECTOR(1 DOWNTO 0);

SIGNAL EX_DATA_FOWARD : STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL EX_REG_DST_MUX : STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL EX_ALU_SRC_A, EX_ALU_SRC_B : STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL EX_ALU_OUT : STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL EX_ALU_OPERATION, EX_ALU_ZERO, EX_ALU_OVERFLOW, EX_ALU_COUT : STD_LOGIC;

-- Sinais do Estagio EX/MEM
SIGNAL EX_ALU_OPERATION : STD_LOGIC;
SIGNAL MEM_DATA_FOWARD : STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL MEM_REG_DST : STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL MEM_WRITE_REG : STD_LOGIC;
SIGNAL MEM_ALU_OUT : STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL MEM_RT_DATA_OUT : STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL MEM_IMED_OUT : STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL MEM_WRITE_OUT, MEM_READ_OUT : STD_LOGIC;
SIGNAL MEM_REG_WRITE : STD_LOGIC;
SIGNAL MEM_MEM_TO_REG : STD_LOGIC_VECTOR(1 DOWNTO 0);

SIGNAL MEM_DATA_OUT : STD_LOGIC_VECTOR(15 DOWNTO 0);

-- Sinais do Estagio MEM/WB
SIGNAL WB_DATA_FOWARD : STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL WB_REG_DST : STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL WB_WRITE_REG : STD_LOGIC;
SIGNAL WB_MEM_OUT : STD_LOGIC_VECTOR(15 DOWNTO 0);

SIGNAL WB_ALU_RESULT : STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL WB_REG_WRITE : STD_LOGIC;
SIGNAL WB_MEM_TO_REG : STD_LOGIC_VECTOR(1 DOWNTO 0);
SIGNAL WB_IMED_OUT : STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL WB_ALU_OUT : STD_LOGIC_VECTOR(15 DOWNTO 0);

BEGIN

	-- Estágio IF
		WITH ID_PC_SOURCE SELECT
			-- Lógica para seleção do próximo PC
			IF_PC_MUX <= 	IF_NEXT_PC 		   WHEN "00", -- PC + 2
							"0000000000000000" WHEN "01", -- Tratamento de erro
							ID_BRANCH_RESULT WHEN "10", -- Branch (a implementar) ---
							ID_JUMP_ADDRESS WHEN "11", -- Jump (a implementar) ---
							"0000000000000000" WHEN OTHERS; -- Default

		IF_PC_INSTANCE: REG PORT MAP(
			D => IF_PC_MUX,
			R_in => PC_WRITE,
			Reset => RESET,
			Clock => CLOCK,
			D_out => IF_PC_CURRENT
		); --OK
		
		IF_PC_ADD_INSTANCE: RIPPLE_CARRY PORT MAP(
			A => IF_PC_CURRENT,
			B => "0000000000000010",
			Cin => '0',
			Add_Sub => '0', -- Operação de soma
			Overflow => IF_PC_ADD_OVERFLOW, -- Salva o resultado do overflow (não utilizado)
			Cout => IF_PC_ADD_COUT, -- Salva o carry out (não utilizado)
			Z => IF_NEXT_PC
		); --OK

		INSTRUCTION_MEMORY_INSTANCE: MEMORY PORT MAP( --NOK
			ADDRESS=>IF_PC_CURRENT,
			DATA_IN=> "0000000000000000", -- Inserção das instruções, nunca acontece 
			DATA_OUT=>IF_INSTRUCTION,
			READ_MEM=>'1', -- Sempre lê
			WRITE_MEM=>'0', -- Nunca escreve
			CLOCK=>CLOCK
		);

		PIPE_IF_ID_INSTANCE: PIPE_IF_ID PORT MAP( --NOK
			-- Inputs
			NEXT_PC_IN => IF_NEXT_PC,
			INSTRUCTION_DATA_IN => IF_INSTRUCTION,

			IF_ID_WRITE => ID_IF_ID_WRITE, --- Vem do controle de hazard
			IF_FLUSH => ID_IF_FLUSH,

			-- Outputs
			NEXT_PC_OUT => ID_NEXT_PC,
			INSTRUCTION_DATA_OUT => ID_INSTRUCTION_DATA,

			-- Controle de clock e reset
			CLOCK => CLOCK,
			RESET => RESET
		);

--===============================================================================
	-- Estagio IF/ID

		ID_RS_OP <= ID_INSTRUCTION_DATA(10 DOWNTO 8); -- Bits de RS
		ID_RT_OP <= ID_INSTRUCTION_DATA(7 DOWNTO 5);  -- Bits de RT
		ID_RD_OP <= ID_INSTRUCTION_DATA(4 DOWNTO 2);  -- Bits de RD


		CONTROL_UNIT_INSTANCE : CONTROL_UNIT PORT MAP( --NOK
			OPCODE => ID_INSTRUCTION_DATA(15 DOWNTO 0),
			REG_EQUAL => ID_REG_EQUAL,

			IF_FLUSH => ID_IF_FLUSH,
			ID_FLUSH => ID_ID_FLUSH,
			EX_FLUSH => ID_EX_FLUSH,
			WB_FLUSH => ID_WB_FLUSH,

			PC_SOURCE => ID_PC_SOURCE,
			ALU_SRC => ID_ALU_SRC,
			REG_DST=> ID_REG_DST,
			ALU_OP=> ID_ALU_OP,

			-- Sinais de controle MEM
			MEM_WRITE=> ID_MEM_WRITE,
			MEM_READ=> ID_MEM_READ,
			-- Sinais de controle WB
			MEM_TO_REG=> ID_MEM_TO_REG,
			REG_WRITE=> ID_REG_WRITE,

		);

		IF_ID_HAZARD_DETECTION_UNIT_INSTANCE : HAZARD_DETECTION_UNIT PORT MAP( --NOK
			-- ID_EX_MEM_READ => , -- EX/MEM ---
			-- ID_EX_RT => , -- EX/MEM ---
			-- IF_ID_RS => , -- IF/ID ---
			-- IF_ID_RT => , -- IF/ID ---
			PC_WRITE => ID_PC_WRITE,
			IF_ID_WRITE => IF_ID_WRITE,
			-- IF_FLUSH => 
		);

		IF_ID_REG_BANK_INSTANCE: REG_BANK PORT MAP( --NOK
			REG_READ1 => ID_RS_OP, -- RS
			REG_READ2 => ID_RT_OP, -- RT
			WRITE_REG => , -- MEM/WB ---
			WRITE_DATA => , -- MEM/WB ---
			REG_WRITE => , -- MEM/WB ---
			DATA_READ1 => ID_REG_DATA1,
			DATA_READ2 => ID_REG_DATA2,
			CLOCK => CLOCK,
			RESET => RESET
		);

		IF_ID_SIGN_EXTEND_INSTANCE: SIGN_EXTEND PORT MAP( --OK
			IN_SIGNAL => ID_INSTRUCTION_DATA(4 DOWNTO 0),
			OUT_SIGNAL => ID_SIGNAL_EXTENDED,
		);

		IF_ID_SHIFT_LEFT_INSTANCE: SHIFT_LEFT2 PORT MAP( --OK
			IN_SIGNAL => ID_SIGNAL_EXTENDED,
			OUT_SIGNAL => ID_SIGNAL_SHIFTED,
		);

		IF_ID_COMPARATOR_INSTANCE: COMPARATOR PORT MAP(
			A => ID_REG_DATA1,
			B => ID_REG_DATA2,
			EQU => ID_REG_EQUAL,
		);

		IF_ID_RIPPLE_BRANCH_INSTANCE: RIPPLE_CARRY PORT MAP( --OK
			A => ID_NEXT_PC,
			B => ID_SIGNAL_SHIFTED,
			Cin => '0',
			Add_Sub => '0',
			Overflow => ID_RIPPLE_BRANCH_OVERFLOW,
			Cout => ID_RIPPLE_BRANCH_COUT,
			Z => ID_BRANCH_RESULT,
		);

		IF_ID_SHIFT_LEFT1_JUMP_INSTANCE: SHIFT_LEFT1 PORT MAP( --OK
			IN_SIGNAL => ID_INSTRUCTION_DATA(12 DOWNTO 0),
			OUT_SIGNAL => ID_JUMP_ADDRESS(13 DOWNTO 0),
		);
		ID_JUMP_ADDRESS(15 DOWNTO 14) <= ID_NEXT_PC(15 DOWNTO 14); -- Concatena os dois bits mais significativos do PC+2

		-- WITH 

		PIPE_ID_EX_INSTANCE: PIPE_ID_EX PORT MAP(
			-- Inputs
			A_IN=> ID_REG_DATA1,
			B_IN=> ID_REG_DATA2,
			SIGNAL_EXT_IN=> ID_SIGNAL_EXTENDED,
			IF_ID_REG_RS_IN=> ID_RS_OP,
			IF_ID_REG_RT_IN=> ID_RT_OP,
			IF_ID_REG_RD_IN=> ID_RD_OP,
			IF_NEXT_PC=> ID_NEXT_PC,

			-- Outputs
			A_OUT=>EX_A,
			B_OUT=>EX_B,
			SIGNAL_EXT_OUT=>EX_SIGNAL_EXTENDED,
			IF_ID_REG_RS_OUT=>EX_RS_OP,
			IF_ID_REG_RT_OUT=>EX_RT_OP,
			IF_ID_REG_RD_OUT=>EX_RD_OP,
			NEXT_PC_OUT=>EX_NEXT_PC,

			-- Sinais de controle EX
			EX_ALU_SRC_IN=>ID_ALU_SRC,
			EX_REG_DST_IN=>ID_REG_DST,
			EX_ALU_OP_IN=>ID_ALU_OP,
			EX_ALU_SRC_OUT=>EX_ALU_SRC,
			EX_REG_DST_OUT=>EX_REG_DST,
			EX_ALU_OP_OUT=>EX_ALU_OP,

			-- Sinais de controle MEM
			MEM_WRITE_IN=>ID_MEM_WRITE,
			MEM_READ_IN=>ID_MEM_READ,
			MEM_WRITE_OUT=>EX_MEM_WRITE,
			MEM_READ_OUT=>EX_MEM_READ,

			-- Sinais de controle WB
			WB_MEM_TO_REG_IN=>ID_MEM_TO_REG,
			WB_REG_WRITE_IN=>ID_REG_WRITE,
			WB_MEM_TO_REG_OUT=>EX_MEM_TO_REG,
			WB_REG_WRITE_OUT=>EX_REG_WRITE,

			CLOCK=> CLOCK
			RESET=> RESET
		);
		
--===============================================================================
--===============================================================================
	-- Estágio ID/EX

		ALU_CONTROL_INSTANCE : ALU_CONTROL PORT MAP(
			ALU_OP => ID_ALU_OP,
			ADD_SUB => ID_SIGNAL_EXTENDED(0), -- ultimo bit do funct
        	ALU_CONTROL_OUT => EX_ALU_OPERATION
		);

		FORWARDING_UNIT_INSTANCE : FORWARDING_UNIT PORT MAP(
			RS => EX_RS_OP,
			RT => EX_RT_OP,
			REG_DST_EX_MEM => MEM_REG_DST, ---
			REG_DST_MEM_WB => WB_REG_DST, ---
			WRITE_REG_EX_MEM => MEM_WRITE_REG, ---
			WRITE_REG_MEM_WB => WB_WRITE_REG, ---
			FOWARD_A => EX_FOWARD_A,
			FOWARD_B => EX_FOWARD_B
		);

		WHEN EX_FOWARD_A SELECT
			EX_ALU_SRC_A <= 	EX_A WHEN "00",
								MEM_DATA_FOWARD WHEN "10",
								WB_DATA_FOWARD WHEN "01",
								EX_A WHEN OTHERS; -- Default

		WHEN EX_FOWARD_B SELECT
			EX_ALU_SRC_B <= 	EX_DATA_FOWARD WHEN "00",
										MEM_DATA_FOWARD WHEN "10",
										WB_DATA_FOWARD WHEN "01",
										EX_DATA_FOWARD WHEN OTHERS; -- Default

		WITH EX_ALU_SRC SELECT
			EX_DATA_FOWARD <= 	EX_SIGNAL_EXTENDED WHEN "1",
								EX_B WHEN "0",
								EX_B WHEN OTHERS; -- Default

		WITH EX_REG_DST SELECT
			EX_REG_DST_MUX <= 	EX_RT_OP WHEN "0",
								EX_RD_OP WHEN "1",
								EX_RT_OP WHEN OTHERS; -- Default

		ALU_INSTANCE : ULA PORT MAP(
			A=> EX_ALU_SRC_A,
			B=> EX_ALU_SRC_B,
			RESULT => EX_ALU_OUT,
			OPERATION=> EX_ALU_OPERATION,
			ZERO => EX_ALU_ZERO,
			OVERFLOW=> EX_ALU_OVERFLOW,
			Cout => EX_ALU_COUT
		);

		PIPE_EX_MEM_INSTANCE: PIPE_EX_MEM PORT MAP(
			-- Inputs
			ALU_OUT_IN=>EX_ALU_OUT,
			RT_DATA_IN=>EX_B,
			IMED_IN=>EX_SIGNAL_EXTENDED,
			REG_DST_IN=>EX_REG_DST_MUX,

			-- Outputs
			ALU_OUT_OUT=> MEM_ALU_OUT,
			RT_DATA_OUT=> MEM_RT_DATA_OUT,
			IMED_OUT=> MEM_IMED_OUT,
			REG_DST_OUT=> MEM_REG_DST,

			-- Sinais de controle
			-- MEM
			MEM_WRITE_IN=> EX_MEM_WRITE,
			MEM_READ_IN=> EX_MEM_READ,
			-- MEM_ALU_RESULT_IN=> ,
			-- MEM_ALU_SRC2_IN=> ,

			MEM_WRITE_OUT=> MEM_WRITE_OUT,
			MEM_READ_OUT=> MEM_READ_OUT,
			-- MEM_ALU_RESULT_OUT=> ,
			-- MEM_ALU_SRC2_OUT=> ,

			-- WB
			WB_MEM_TO_REG_IN=> EX_MEM_TO_REG,
			WB_REG_WRITE_IN=> EX_REG_WRITE,

			WB_MEM_TO_REG_OUT=> MEM_MEM_TO_REG,
			WB_REG_WRITE_OUT=> MEM_REG_WRITE,

			-- Controle de clock e reset
			CLOCK=> CLOCK,
			RESET=> RESET,
		)
		
--===============================================================================
--===============================================================================
	-- Estagio EX/MEM

		DATA_MEMORY_INSTANCE: MEMORY PORT MAP( --NOK
			ADDRESS=> MEM_ALU_OUT,
			DATA_IN=> MEM_RT_DATA_OUT,
			DATA_OUT=> MEM_DATA_OUT,
			READ_MEM=> MEM_READ_OUT, 
			WRITE_MEM=> MEM_WRITE_OUT, 
			CLOCK=>CLOCK
		);

		PIPE_MEM_WB_INSTANCE : PIPE_MEM_WB PORT MAP(
			-- Inputs
			MEM_OUT_IN => MEM_DATA_OUT,
			ALU_RESULT_IN => MEM_ALU_OUT,
			IMED_IN => MEM_IMED_OUT,
			REG_DST_IN => MEM_REG_DST,
			
			-- Outputs
			MEM_OUT_OUT => WB_MEM_OUT,
			ALU_RESULT_OUT => WB_ALU_OUT,
			IMED_OUT => WB_IMED_OUT,
			REG_DST_OUT => WB_REG_DST,

			-- Sinais de controle
			-- WB
			WB_MEM_TO_REG_IN => MEM_MEM_TO_REG,
			WB_REG_WRITE_IN => MEM_REG_WRITE,

			WB_MEM_TO_REG_OUT => WB_MEM_TO_REG,
			WB_REG_WRITE_OUT => WB_REG_WRITE,

			CLOCK => CLOCK,
			RESET => RESET,
		);

	-- Estagio MEM/WB

		WITH WB_MEM_TO_REG_OUT SELECT
			WB_MEM_TO_REG <= 	WB_MEM_OUT WHEN  "00",
								WB_IMED_OUT WHEN "01",
								WB_ALU_OUT WHEN "10",
								WB_ALU_OUT WHEN OTHERS; -- Default

	-- PROCESSOS PARA O DIVISOR DE CLOCK
    ClockDivide: PROCESS
            BEGIN
            WAIT UNTIL CLOCK_50'EVENT and CLOCK_50 = '1'; -- Na subida do clock,
            IF clockticks < max THEN
                clockticks <= clockticks + 1; -- Soma o contador clockticks até o máximo estipulado pelo usuário
            ELSE
                clockticks <= 0;					-- Quando chega no máximo zera
            END IF;
            IF clockticks < half THEN			-- Half representa a metade do ciclo, quando chega liga o clock
                CLOCK <= '0';
            ELSE
                CLOCK <= '1';
            END IF;
        END PROCESS;
		  
-- Basicamente, o ClockDivide é um processo que conta até um certo número e altera o valor do clock com base na
-- metade desse número, criando um efeito parecido com isso:
--
-- Para max = 4
-- CLK_50 - -: _|¯|_|¯|_|¯|_|¯|_|¯|_|¯|...
--	CLK- - - -: ___|¯¯¯|___|¯¯¯|___|¯¯¯|...
---          -------------t--------------
-- Com isso, quanto maior for "max", maior será o ciclo de CLK
END Behavior;
