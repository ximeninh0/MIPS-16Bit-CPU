LIBRARY ieee;
USE ieee.std_logic_1164.all;
use work.CPU_PACKAGE.all;

ENTITY TWO_DIGITS_7_SEGS IS 
		port(
			NUMBER : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
			TRANSLATED_FIRST_DIGIT: OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
			TRANSLATED_SECOND_DIGIT: OUT STD_LOGIC_VECTOR(6 DOWNTO 0)

		);
END TWO_DIGITS_7_SEGS;

ARCHITECTURE Behavior OF TWO_DIGITS_7_SEGS IS
-- Decodificador de numeros de 4 bits para 7 segmentos

BEGIN
	WITH NUMBER SELECT
    TRANSLATED_FIRST_DIGIT <=
        "0000001" when "0000000000000000", --0
        "0000001" when "0000000000000001", --1
        "0000001" when "0000000000000010", --2
        "0000001" when "0000000000000011", --3
        "0000001" when "0000000000000100", --4
        "0000001" when "0000000000000101", --5
        "0000001" when "0000000000000110", --6
        "0000001" when "0000000000000111", --7
        "0000001" when "0000000000001000", --8
        "0000001" when "0000000000001001", --9
		  
        "1001111" when "0000000000001010", -- 10
        "1001111" when "0000000000001011", -- 11
        "1001111" when "0000000000001100", -- 12
        "1001111" when "0000000000001101", -- 13
        "1001111" when "0000000000001110", -- 14
        "1001111" when "0000000000001111", -- 15
        "1001111" when "0000000000010000", -- 16
        "1001111" when "0000000000010001", -- 17
        "1001111" when "0000000000010010", -- 18
        "1001111" when "0000000000010011", -- 19
		  
        "0010010" when "0000000000010100", -- 20
        "0010010" when "0000000000010101", -- 21
        "0010010" when "0000000000010110", -- 22
        "0010010" when "0000000000010111", -- 23
        "0010010" when "0000000000011000", -- 24
        "0010010" when "0000000000011001", -- 25
        "0010010" when "0000000000011010", -- 26
        "0010010" when "0000000000011011", -- 27
        "0010010" when "0000000000011100", -- 28
        "0010010" when "0000000000011101", -- 29
		  
        "0000110" when "0000000000011110", -- 30
        "0000110" when "0000000000011111", -- 31
        "0000110" when "0000000000100000", -- 32
        "0000110" when "0000000000100001", -- 33
        "0000110" when "0000000000100010", -- 34
        "0000110" when "0000000000100011", -- 35
        "0000110" when "0000000000100100", -- 36
        "0000110" when "0000000000100101", -- 37
        "0000110" when "0000000000100110", -- 38
        "0000110" when "0000000000100111", -- 39
		  
        "1001100" when "0000000000101000", -- 40
        "1001100" when "0000000000101001", -- 41
        "1001100" when "0000000000101010", -- 42
        "1001100" when "0000000000101011", -- 43
        "1001100" when "0000000000101100", -- 44
        "1001100" when "0000000000101101", -- 45
        "1001100" when "0000000000101110", -- 46
        "1001100" when "0000000000101111", -- 47
        "1001100" when "0000000000110000", -- 48
        "1001100" when "0000000000110001", -- 49
		  
        "0100100" when "0000000000110010", -- 50
        "0100100" when "0000000000110011", -- 51
        "0100100" when "0000000000110100", -- 52
        "0100100" when "0000000000110101", -- 53
        "0100100" when "0000000000110110", -- 54
        "0100100" when "0000000000110111", -- 55
        "0100100" when "0000000000111000", -- 56
        "0100100" when "0000000000111001", -- 57
        "0100100" when "0000000000111010", -- 58
        "0100100" when "0000000000111011", -- 59
		  
        "0100000" when "0000000000111100", -- 60
        "0100000" when "0000000000111101", -- 61
        "0100000" when "0000000000111110", -- 62
        "0100000" when "0000000000111111", -- 63
        "0100000" when "0000000001000000", -- 64
        "0100000" when "0000000001000001", -- 65
        "0100000" when "0000000001000010", -- 66
        "0100000" when "0000000001000011", -- 67
        "0100000" when "0000000001000100", -- 68
        "0100000" when "0000000001000101", -- 69
		  
        "0001111" when "0000000001000110", -- 70
        "0001111" when "0000000001000111", -- 71
        "0001111" when "0000000001001000", -- 72
        "0001111" when "0000000001001001", -- 73
        "0001111" when "0000000001001010", -- 74
        "0001111" when "0000000001001011", -- 75
        "0001111" when "0000000001001100", -- 76
        "0001111" when "0000000001001101", -- 77
        "0001111" when "0000000001001110", -- 78
        "0001111" when "0000000001001111", -- 79
		  
        "0000000" when "0000000001010000", -- 80
        "0000000" when "0000000001010001", -- 81
        "0000000" when "0000000001010010", -- 82
        "0000000" when "0000000001010011", -- 83
        "0000000" when "0000000001010100", -- 84
        "0000000" when "0000000001010101", -- 85
        "0000000" when "0000000001010110", -- 86
        "0000000" when "0000000001010111", -- 87
        "0000000" when "0000000001011000", -- 88
        "0000000" when "0000000001011001", -- 89
		  
        "0000100" when "0000000001011010", -- 90
        "0000100" when "0000000001011011", -- 91
        "0000100" when "0000000001011100", -- 92
        "0000100" when "0000000001011101", -- 93
        "0000100" when "0000000001011110", -- 94
        "0000100" when "0000000001011111", -- 95
        "0000100" when "0000000001100000", -- 96
        "0000100" when "0000000001100001", -- 97
        "0000100" when "0000000001100010", -- 98
        "0000100" when "0000000001100011", -- 99

        "1111111" when others; -- apagado
		  
		  
-- Para o segundo dígito (de 0 a 9)
WITH NUMBER SELECT
    TRANSLATED_SECOND_DIGIT <=
        "0000001" when "0000000000000000", -- 0
        "1001111" when "0000000000000001", -- 1
        "0010010" when "0000000000000010", -- 2
        "0000110" when "0000000000000011", -- 3
        "1001100" when "0000000000000100", -- 4
        "0100100" when "0000000000000101", -- 5
        "0100000" when "0000000000000110", -- 6
        "0001111" when "0000000000000111", -- 7
        "0000000" when "0000000000001000", -- 8
        "0000100" when "0000000000001001", -- 9
		  
        "0000001" when "0000000000001010", -- 10
        "1001111" when "0000000000001011", -- 11
        "0010010" when "0000000000001100", -- 12
        "0000110" when "0000000000001101", -- 13
        "1001100" when "0000000000001110", -- 14
        "0100100" when "0000000000001111", -- 15
        "0100000" when "0000000000010000", -- 16
        "0001111" when "0000000000010001", -- 17
        "0000000" when "0000000000010010", -- 18
        "0000100" when "0000000000010011", -- 19
		  
        "0000001" when "0000000000010100", -- 20
        "1001111" when "0000000000010101", -- 21
        "0010010" when "0000000000010110", -- 22
        "0000110" when "0000000000010111", -- 23
        "1001100" when "0000000000011000", -- 24
        "0100100" when "0000000000011001", -- 25
        "0100000" when "0000000000011010", -- 26
        "0001111" when "0000000000011011", -- 27
        "0000000" when "0000000000011100", -- 28
        "0000100" when "0000000000011101", -- 29
		  
        "0000001" when "0000000000011110", -- 30
        "1001111" when "0000000000011111", -- 31
        "0010010" when "0000000000100000", -- 32
        "0000110" when "0000000000100001", -- 33
        "1001100" when "0000000000100010", -- 34
        "0100100" when "0000000000100011", -- 35
        "0100000" when "0000000000100100", -- 36
        "0001111" when "0000000000100101", -- 37
        "0000000" when "0000000000100110", -- 38
        "0000100" when "0000000000100111", -- 39
		  
        "0000001" when "0000000000101000", -- 40
        "1001111" when "0000000000101001", -- 41
        "0010010" when "0000000000101010", -- 42
        "0000110" when "0000000000101011", -- 43
        "1001100" when "0000000000101100", -- 44
        "0100100" when "0000000000101101", -- 45
        "0100000" when "0000000000101110", -- 46
        "0001111" when "0000000000101111", -- 47
        "0000000" when "0000000000110000", -- 48
        "0000100" when "0000000000110001", -- 49
		  
        "0000001" when "0000000000110010", -- 50
        "1001111" when "0000000000110011", -- 51
        "0010010" when "0000000000110100", -- 52
        "0000110" when "0000000000110101", -- 53
        "1001100" when "0000000000110110", -- 54
        "0100100" when "0000000000110111", -- 55
        "0100000" when "0000000000111000", -- 56
        "0001111" when "0000000000111001", -- 57
        "0000000" when "0000000000111010", -- 58
        "0000100" when "0000000000111011", -- 59
		  
        "0000001" when "0000000000111100", -- 60
        "1001111" when "0000000000111101", -- 61
        "0010010" when "0000000000111110", -- 62
        "0000110" when "0000000000111111", -- 63
        "1001100" when "0000000001000000", -- 64
        "0100100" when "0000000001000001", -- 65
        "0100000" when "0000000001000010", -- 66
        "0001111" when "0000000001000011", -- 67
        "0000000" when "0000000001000100", -- 68
        "0000100" when "0000000001000101", -- 69
		  
        "0000001" when "0000000001000110", -- 70
        "1001111" when "0000000001000111", -- 71
        "0010010" when "0000000001001000", -- 72
        "0000110" when "0000000001001001", -- 73
        "1001100" when "0000000001001010", -- 74
        "0100100" when "0000000001001011", -- 75
        "0100000" when "0000000001001100", -- 76
        "0001111" when "0000000001001101", -- 77
        "0000000" when "0000000001001110", -- 78
        "0000100" when "0000000001001111", -- 79
		  
        "0000001" when "0000000001010000", -- 80
        "1001111" when "0000000001010001", -- 81
        "0010010" when "0000000001010010", -- 82
        "0000110" when "0000000001010011", -- 83
        "1001100" when "0000000001010100", -- 84
        "0100100" when "0000000001010101", -- 85
        "0100000" when "0000000001010110", -- 86
        "0001111" when "0000000001010111", -- 87
        "0000000" when "0000000001011000", -- 88
        "0000100" when "0000000001011001", -- 89
		  
        "0000001" when "0000000001011010", -- 90
        "1001111" when "0000000001011011", -- 91
        "0010010" when "0000000001011100", -- 92
        "0000110" when "0000000001011101", -- 93
        "1001100" when "0000000001011110", -- 94
        "0100100" when "0000000001011111", -- 95
        "0100000" when "0000000001100000", -- 96
        "0001111" when "0000000001100001", -- 97
        "0000000" when "0000000001100010", -- 98
        "0000100" when "0000000001100011", -- 99
        "1111111" when others; -- apagado


END Behavior;