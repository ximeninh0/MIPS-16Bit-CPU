LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY PIPE_IF_ID IS 
    port(
        NEXT_PC_IN : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
        INSTRUCTION_DATA_IN : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
        IF_D_WRITE : IN STD_LOGIC;
        IF_FLUSH : IN STD_LOGIC;
        NEXT_PC_OUT : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
        INSTRUCTION_DATA_OUT : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
    );
END PIPE_IF_ID;


ARCHITECTURE Behavior OF PIPE_IF_ID IS

BEGIN
END Behavior;
