LIBRARY ieee;
USE ieee.std_logic_1164.all;
use work.CPU_PACKAGE.all;

ENTITY TWO_DIGITS_7_SEGS IS 
		port(
			NUMBER : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
			TRANSLATED_FIRST_DIGIT: OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
			TRANSLATED_SECOND_DIGIT: OUT STD_LOGIC_VECTOR(6 DOWNTO 0)

		);
END TWO_DIGITS_7_SEGS;

ARCHITECTURE Behavior OF TWO_DIGITS_7_SEGS IS
-- Decodificador de numeros de 4 bits para 7 segmentos

BEGIN
	WITH NUMBER SELECT
    TRANSLATED_FIRST_DIGIT <=
        "0000001" when "0000000000000000", --0
        "0000001" when "0000000000000001", --1
        "0000001" when "0000000000000010", --2
        "0000001" when "0000000000000011", --3
        "0000001" when "0000000000000100", --4
        "0000001" when "0000000000000101", --5
        "0000001" when "0000000000000110", --6
        "0000001" when "0000000000000111", --7
        "0000001" when "0000000000001000", --8
        "0000001" when "0000000000001001", --9
		  
        "1001111" when "0000000000001010", --10
        "1001111" when "0000000000001011", --11
        "1001111" when "0000000000001100", --12
        "1001111" when "0000000000001101", --13
        "1001111" when "0000000000001110", --14
        "1001111" when "0000000000001111", --15
        "1001111" when "0000000000010000", --16
        "1001111" when "0000000000010001", --17
        "1001111" when "0000000000010010", --18
        "1001111" when "0000000000010011", --19
		  
        "0010010" when "0000000000010100", --20
        "0010010" when "0000000000010101", --21
        "0010010" when "0000000000010110", --22
        "0010010" when "0000000000010111", --23
        "0010010" when "0000000000011000", --24
        "0010010" when "0000000000011001", --25
        "0010010" when "0000000000011010", --26
        "0010010" when "0000000000011011", --27
        "0010010" when "0000000000011100", --28
        "0010010" when "0000000000011101", --29
--		  
--        "0000001" when "0000000000011110", --0
--        "1001111" when "0000000000000001", --1
--        "0010010" when "0000000000000010", --2
--        "0000110" when "0000000000000011", --3
--        "1001100" when "0000000000000100", --4
--        "0100100" when "0000000000000101", --5
--        "0100000" when "0000000000000110", --6
--        "0001111" when "0000000000000111", --7
--        "0000000" when "0000000000001000", --8
--        "0000100" when "0000000000001001", --9

        "1111111" when others; -- apagado
		  
		  
	WITH NUMBER SELECT
    TRANSLATED_SECOND_DIGIT <=
        "0000001" when "0000000000000000", --0
        "1001111" when "0000000000000001", --1
        "0010010" when "0000000000000010", --2
        "0000110" when "0000000000000011", --3
        "1001100" when "0000000000000100", --4
        "0100100" when "0000000000000101", --5
        "0100000" when "0000000000000110", --6
        "0001111" when "0000000000000111", --7
        "0000000" when "0000000000001000", --8
        "0000100" when "0000000000001001", --9
		  
        "0000001" when "0000000000001010", --10
        "1001111" when "0000000000001011", --11
        "0010010" when "0000000000001100", --12
        "0000110" when "0000000000001101", --13
        "1001100" when "0000000000001110", --14
        "0100100" when "0000000000001111", --15
        "0100000" when "0000000000010000", --16
        "0001111" when "0000000000010001", --17
        "0000000" when "0000000000010010", --18
        "0000100" when "0000000000010011", --19
		  
        "0000001" when "0000000000010100", --20
        "1001111" when "0000000000010101", --21
        "0010010" when "0000000000010110", --22
        "0000110" when "0000000000010111", --23
        "1001100" when "0000000000011000", --24
        "0100100" when "0000000000011001", --25
        "0100000" when "0000000000011010", --26
        "0001111" when "0000000000011011", --27
        "0000000" when "0000000000011100", --28
        "0000100" when "0000000000011101", --29
        "1111111" when others; -- apagado

END Behavior;