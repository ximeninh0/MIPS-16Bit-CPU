LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY PIPE_MEM_WB IS 

port(
    -- Inputs
    MEM_OUT_IN : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    ALU_RESULT_IN : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    REG_DST_IN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);

    -- Outputs
    MEM_OUT_OUT : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
    ALU_RESULT_OUT : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
    REG_DST_OUT : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);

    -- Sinais de controle
    -- WB
    WB_MEM_TO_REG_IN : IN STD_LOGIC;
    WB_REG_WRITE_IN : IN STD_LOGIC;

    WB_MEM_TO_REG_OUT : OUT STD_LOGIC;
    WB_REG_WRITE_OUT : OUT STD_LOGIC;

    -- Controle de clock e reset
    CLOCK : IN STD_LOGIC;
    RESET : IN STD_LOGIC
);
END PIPE_MEM_WB;

ARCHITECTURE Behavior OF PIPE_MEM_WB IS

    -- Dados
    MEM_OUT_INSTANCE: REG PORT MAP(MEM_OUT_IN,'1',RESET,CLOCK,MEM_OUT_OUT);
    ALU_RESULT_INSTANCE: REG PORT MAP(ALU_RESULT_IN,'1',RESET,CLOCK,ALU_RESULT_OUT);
    REG_DST_INSTANCE: FOUR_BIT_REG PORT MAP(REG_DST_IN,'1',RESET,CLOCK,REG_DST_OUT);

    -- WB
    WB_MEM_TO_REG_INSTANCE: ONE_BIT_REG PORT MAP(WB_MEM_TO_REG_IN,'1',RESET,CLOCK,WB_MEM_TO_REG_OUT);
    WB_REG_WRITE_INSTANCE: ONE_BIT_REG PORT MAP(WB_REG_WRITE_IN,'1',RESET,CLOCK,WB_REG_WRITE_OUT);

BEGIN
END Behavior;
