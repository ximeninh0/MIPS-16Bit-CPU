LIBRARY ieee;
use ieee.std_logic_1164.all;

PACKAGE CPU_PACKAGE IS

constant WORD_SIZE     : integer := 16;
constant ADDR_SIZE     : integer := 16;
constant BYTE_SIZE     : integer := 8;

END CPU_PACKAGE;
