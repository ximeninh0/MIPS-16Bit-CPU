LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY PIPE_EX_MEM IS 

END PIPE_EX_MEM;
    port(
        -- Inputs
        ALU_OUT_IN : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
        RT_DATA_IN : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
        IMED_IN : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
        REG_DST_IN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);

        -- Outputs
        ALU_OUT_OUT : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);    
        RT_DATA_OUT : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
        IMED_OUT : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
        REG_DST_OUT : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);

        -- Sinais de controle
        -- MEM
        MEM_WRITE_IN : IN STD_LOGIC;
        MEM_READ_IN : IN STD_LOGIC;
        -- MEM_ALU_RESULT_IN : IN STD_LOGIC;
        -- MEM_ALU_SRC2_IN : IN STD_LOGIC;

        MEM_WRITE_OUT : OUT STD_LOGIC;
        MEM_READ_OUT : OUT STD_LOGIC;
        -- MEM_ALU_RESULT_OUT : OUT STD_LOGIC;
        -- MEM_ALU_SRC2_OUT : OUT STD_LOGIC;

        -- WB
        WB_MEM_TO_REG_IN : IN STD_LOGIC_VECTOR(1 DOWNTO 0);;
        WB_REG_WRITE_IN : IN STD_LOGIC;

        WB_MEM_TO_REG_OUT : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);;
        WB_REG_WRITE_OUT : OUT STD_LOGIC;

        -- Controle de clock e reset
        CLOCK : IN STD_LOGIC;
        RESET : IN STD_LOGIC
    );

ARCHITECTURE Behavior OF PIPE_EX_MEM IS

BEGIN
    -- Dados
    ALU_OUT_INSTANCE: REG PORT MAP(ALU_OUT_IN,'1',RESET,CLOCK,ALU_OUT_OUT);
    RT_DATA_INSTANCE: REG PORT MAP(RT_DATA_IN,'1',RESET,CLOCK,RT_DATA_OUT);
    IMED_INSTANCE: REG PORT MAP(IMED_IN,'1',RESET,CLOCK,IMED_OUT);
    REG_DST_INSTANCE: FOUR_BIT_REG PORT MAP(REG_DST_IN,'1',RESET,CLOCK,REG_DST_OUT);

    -- MEM
    MEM_WRITE_INSTANCE: ONE_BIT_REG PORT MAP(MEM_WRITE_IN,'1',RESET,CLOCK,MEM_WRITE_OUT);
    MEM_READ_INSTANCE: ONE_BIT_REG PORT MAP(MEM_READ_IN,'1',RESET,CLOCK,MEM_READ_OUT);
    -- MEM_ALU_RESULT_INSTANCE: ONE_BIT_REG PORT MAP(MEM_ALU_RESULT_IN,'1',RESET,CLOCK,MEM_ALU_RESULT_OUT);
    -- MEM_ALU_SRC2_INSTANCE: ONE_BIT_REG PORT MAP(MEM_ALU_SRC2_IN,'1',RESET,CLOCK,MEM_ALU_SRC2_OUT);

    -- WB
    WB_MEM_TO_REG_INSTANCE: TWO_BIT_REG PORT MAP(WB_MEM_TO_REG_IN,'1',RESET,CLOCK,WB_MEM_TO_REG_OUT);
    WB_REG_WRITE_INSTANCE: ONE_BIT_REG PORT MAP(WB_REG_WRITE_IN,'1',RESET,CLOCK,WB_REG_WRITE_OUT);

END Behavior;
