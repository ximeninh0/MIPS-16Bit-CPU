LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY PIPE_MEM_WB IS 

port(
    MEM_OUT_IN : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    ALU_OUT_IN : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    REG_DST_IN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);

    MEM_OUT_OUT : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
    ALU_OUT_OUT : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
    REG_DST_OUT : OUT STD_LOGIC_VECTOR(3 DOWNTO 0) 
);
END PIPE_MEM_WB;

ARCHITECTURE Behavior OF PIPE_MEM_WB IS

BEGIN
END Behavior;
