LIBRARY ieee;
use ieee.std_logic_1164.all;
--PACKAGE COM TODOS OS COMPONENTES UTILIZADOS NA CPU E NA ULA

PACKAGE CPU_PACKAGE IS
	COMPONENT ULA IS 
		port(
			A,B : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			OPERATION: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
			ZERO, OVERFLOW,Cout : OUT STD_LOGIC;
			RESULT: OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
			Equ,Grt,Lst : OUT STD_LOGIC
		);
	END COMPONENT;
	
	COMPONENT UC_CPU IS 
		port(
			OPCODE : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			Clock : in std_logic;
			RESET : IN STD_LOGIC;
			En : IN STD_LOGIC;
			R_in : OUT STD_LOGIC_VECTOR(1 TO 3);
			R_out : OUT STD_LOGIC_VECTOR(1 TO 3);
			G_in : OUT STD_LOGIC;
			G_out : OUT STD_LOGIC;
			A_in : OUT STD_LOGIC;
			B_in : OUT STD_LOGIC;
			DONE : OUT STD_LOGIC;
			EXTERN : OUT STD_LOGIC;
			OP_ULA: OUT STD_LOGIC_VECTOR (3 DOWNTO 0)
		);
	END COMPONENT;
	
	COMPONENT UC_LCD IS 
		  port(
			OPCODE : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			 CLOCK : IN STD_LOGIC;
			 EQU,GRT,LST,ENABLE : IN STD_LOGIC;
			 LCD_DATA : out STD_LOGIC_VECTOR(7 DOWNTO 0);
			 LCD_RW : OUT STD_LOGIC;
			 LCD_EN : OUT STD_LOGIC;
			 LCD_RS: OUT STD_LOGIC
		  );
	END COMPONENT;
	
	COMPONENT REG_BANK IS 
		port(
				REG_READ1,REG_READ2 :IN STD_LOGIC_VECTOR(1 DOWNTO 0);
				WRITE_REG :IN STD_LOGIC_VECTOR(1 DOWNTO 0);
				WRITE_DATA :IN STD_LOGIC_VECTOR(3 DOWNTO 0);
				REG_WRITE,REG_READ: IN STD_LOGIC;
				DATA_READ1 :OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
				DATA_READ2 :OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
		);
	END COMPONENT;
	
	COMPONENT AND_COMPONENT IS 
		port(
			X,Y :IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			Z : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
		);
	END COMPONENT;
	
	COMPONENT OR_COMPONENT IS
		port(
			X,Y :IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			Z : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
		);
	END COMPONENT;
	
	COMPONENT NOT_COMPONENT IS
		port(
			X,Y :IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			Z : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
		);
	END COMPONENT;
	
	COMPONENT MULTI_COMPONENT IS
		port(
			X,Y :IN STD_LOGIC_VECTOR(1 DOWNTO 0);
			Z : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
		);
	END COMPONENT;
	
	
	COMPONENT RIPPLE_CARRY IS 
		port(
			A,B : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			Cin : IN STD_LOGIC;
			Add_sub: IN STD_LOGIC;
			Overflow: OUT STD_LOGIC;
			Cout : OUT STD_LOGIC;
			Z : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
		);
	END COMPONENT;
	
	COMPONENT FULLADDER IS 
		port(
			A,B,Cin : IN STD_LOGIC;
			S,Cout : OUT STD_LOGIC
		);
	END COMPONENT;
	
	COMPONENT COMPARATOR IS 
		port(
			A,B : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			EQU,GRT,LST : OUT STD_LOGIC
		);
	END COMPONENT;
	
	COMPONENT SEGS_3_TRANSLATOR IS
		port(
			NUMBER : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
			TRANSLATED : OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
		);
	END COMPONENT;
	
	COMPONENT SEGS_4_TRANSLATOR IS 
		port(
			NUMBER : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			TRANSLATED : OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
		);
	END COMPONENT;
	
	COMPONENT MUX_2_TO_1 IS 
		port(
			KEY : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
			X1,X2 : IN STD_LOGIC;
			F : OUT STD_LOGIC
		);
	END COMPONENT;
	
	COMPONENT MUX_5_TO_1 IS 
		port(
			KEY : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
			X1,X2,X3,X4,X5 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			F : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
		);
	END COMPONENT;
	
	COMPONENT BUFFER_TRI IS 
		port(
			ENTRADA : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			GATE : IN STD_LOGIC;
			SAIDA: OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
		);
	END COMPONENT;
	
	COMPONENT REG IS 
		port(
			D : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			R_in,Reset,Clock : IN STD_LOGIC;
			D_out: OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
		);
	END COMPONENT;
	
END CPU_PACKAGE;
