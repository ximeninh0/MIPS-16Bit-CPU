LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY PIPE_ID_EX IS 
    port(
        A_IN : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
        B_IN : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
        SIGNAL_EXT_IN : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
        IF_ID_REG_RS_IN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
        IF_ID_REG_RT_1_IN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
        IF_ID_REG_RT_2_IN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
        IF_ID_REG_RS_IN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);

        A_OUT : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
        B_OUT : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
        SIGNAL_EXT_OUT : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
        IF_ID_REG_RS_OUT : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
        IF_ID_REG_RT_1_OUT : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
        IF_ID_REG_RT_2_OUT : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
        IF_ID_REG_RS_OUT : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)

        EX_ALU_SRC_IN : IN STD_LOGIC;
        EX_REG_DST_IN : IN STD_LOGIC;
        EX_ALU_OP_IN : IN STD_LOGIC_VECTOR(1 DOWNTO 0);

        MEM_WRITE_IN : IN STD_LOGIC;
        MEM_READ_IN : IN STD_LOGIC;
        MEM_ALU_IN : IN STD_LOGIC;
        MEM_ALU_SRC2_IN : IN STD_LOGIC;

        WB_ALU_SRC_IN : IN STD_LOGIC;
        WB_ALU_SRC_IN : IN STD_LOGIC;

    );
END PIPE_ID_EX;


ARCHITECTURE Behavior OF PIPE_ID_EX IS

BEGIN
END Behavior;
